* Extracted by KLayout on : 19/02/2025 20:30

.SUBCKT alu
X$1 NWELL VIA_via9_10_1600_1600_1_1_3360_3360
X$2 NWELL VIA_via9_10_1600_1600_1_1_3360_3360
X$3 NWELL VIA_via9_10_1600_1600_1_1_3360_3360
X$4 NWELL VIA_via9_10_1600_1600_1_1_3360_3360
X$5 b[0] \$3 NWELL \$224 PWELL BUF_X1
X$6 \$224 \$3 NWELL \$496 PWELL BUF_X1
X$7 \$496 NWELL \$90 \$3 PWELL BUF_X4
X$8 \$533 \$279 \$3 NWELL \$278 PWELL NOR2_X1
X$9 a[3] \$3 NWELL \$352 PWELL INV_X1
X$10 \$3 NWELL PWELL FILLCELL_X1
X$11 a[3] \$3 NWELL \$397 PWELL CLKBUF_X1
X$12 \$284 \$3 NWELL \$174 PWELL BUF_X2
X$13 b[1] \$3 NWELL \$284 PWELL CLKBUF_X2
X$14 \$661 NWELL \$173 \$3 PWELL BUF_X4
X$15 \$174 \$351 \$416 NWELL \$586 \$3 PWELL OAI21_X1
X$16 \$3 NWELL PWELL FILLCELL_X4
X$17 \$3 NWELL PWELL FILLCELL_X2
X$18 \$3 NWELL PWELL FILLCELL_X4
X$19 \$3 NWELL PWELL NWELL TAPCELL_X1
X$20 \$3 NWELL PWELL FILLCELL_X2
X$21 \$3 NWELL PWELL NWELL TAPCELL_X1
X$22 \$3 NWELL PWELL FILLCELL_X8
X$23 \$3 NWELL PWELL FILLCELL_X1
X$24 a[3] \$90 a[2] \$3 NWELL \$533 PWELL MUX2_X1
X$25 NWELL VIA_via1_2_940_340_1_3_300_300
X$26 NWELL VIA_via2_3_940_340_1_3_320_320
X$27 NWELL VIA_via3_4_940_340_1_3_320_320
X$28 \$3 NWELL PWELL FILLCELL_X2
X$29 \$382 \$534 \$3 NWELL \$574 PWELL NOR2_X1
X$30 \$533 \$279 \$3 NWELL \$645 PWELL NAND2_X1
X$31 \$3 NWELL PWELL FILLCELL_X8
X$32 \$3 NWELL PWELL FILLCELL_X1
X$33 \$174 \$3 NWELL \$661 PWELL BUF_X2
X$34 \$3 NWELL PWELL FILLCELL_X4
X$35 \$126 \$173 \$3 NWELL \$612 PWELL NAND2_X1
X$36 \$3 NWELL PWELL FILLCELL_X1
X$37 a[7] \$3 NWELL \$222 PWELL CLKBUF_X1
X$38 b[7] \$3 NWELL \$554 PWELL CLKBUF_X1
X$39 \$126 \$284 \$3 NWELL \$614 PWELL NOR2_X1
X$40 \$197 \$200 \$3 NWELL \$471 PWELL NAND2_X1
X$41 \$3 NWELL PWELL FILLCELL_X1
X$42 \$3 NWELL PWELL FILLCELL_X4
X$43 \$3 NWELL PWELL FILLCELL_X1
X$44 \$357 \$356 \$471 \$174 \$3 \$421 NWELL PWELL AOI211_X1
X$45 \$3 NWELL PWELL FILLCELL_X8
X$46 \$3 NWELL PWELL FILLCELL_X2
X$47 \$3 NWELL PWELL FILLCELL_X2
X$48 \$3 NWELL PWELL FILLCELL_X1
X$49 \$174 \$289 \$614 \$357 \$3 \$683 NWELL PWELL AOI211_X1
X$50 \$3 NWELL PWELL FILLCELL_X2
X$51 \$3 NWELL PWELL FILLCELL_X1
X$52 \$471 \$770 \$174 \$3 NWELL \$698 PWELL NOR3_X1
X$53 NWELL VIA_via1_2_940_340_1_3_300_300
X$54 NWELL VIA_via2_3_940_340_1_3_320_320
X$55 NWELL VIA_via3_4_940_340_1_3_320_320
X$56 \$683 \$811 \$231 \$3 \$362 NWELL PWELL AOI21_X1
X$57 \$3 NWELL PWELL FILLCELL_X4
X$58 \$3 NWELL PWELL FILLCELL_X2
X$59 \$3 NWELL PWELL NWELL TAPCELL_X1
X$60 \$3 NWELL PWELL FILLCELL_X2
X$61 \$3 NWELL PWELL FILLCELL_X1
X$62 \$3 NWELL PWELL FILLCELL_X1
X$63 \$421 \$220 \$585 \$3 NWELL \$595 PWELL OR3_X1
X$64 \$474 \$231 NWELL \$3 \$523 PWELL AND2_X1
X$65 \$3 NWELL PWELL FILLCELL_X2
X$66 \$255 \$474 \$698 \$545 \$335 \$3 NWELL \$705 PWELL AOI221_X1
X$67 \$3 NWELL PWELL FILLCELL_X1
X$68 \$458 \$3 NWELL \$545 PWELL BUF_X2
X$69 \$708 \$705 \$586 \$3 NWELL \$593 PWELL NAND3_X1
X$70 b[3] \$397 \$3 NWELL \$619 PWELL NOR2_X2
X$71 \$595 \$523 \$233 \$552 \$511 NWELL \$3 PWELL AOI211_X2
X$72 \$324 \$3 NWELL \$439 PWELL CLKBUF_X1
X$73 \$3 NWELL PWELL FILLCELL_X2
X$74 \$711 \$176 \$549 \$233 \$3 NWELL \$709 PWELL AOI22_X1
X$75 \$620 \$545 \$549 \$3 NWELL PWELL NOR2_X4
X$76 \$545 \$551 \$549 \$3 \$313 NWELL PWELL AOI21_X1
X$77 \$365 \$3 NWELL \$291 PWELL CLKBUF_X1
X$78 \$3 NWELL PWELL FILLCELL_X1
X$79 \$3 NWELL PWELL FILLCELL_X2
X$80 \$3 NWELL PWELL FILLCELL_X8
X$81 \$448 \$3 NWELL \$509 PWELL CLKBUF_X1
X$82 \$3 NWELL PWELL FILLCELL_X1
X$83 \$3 NWELL PWELL FILLCELL_X4
X$84 \$3 NWELL PWELL FILLCELL_X2
X$85 NWELL VIA_via1_2_940_340_1_3_300_300
X$86 NWELL VIA_via2_3_940_340_1_3_320_320
X$87 NWELL VIA_via3_4_940_340_1_3_320_320
X$88 \$733 \$366 \$732 NWELL \$585 \$3 PWELL OAI21_X1
X$89 \$554 \$197 \$3 NWELL \$733 PWELL NAND2_X1
X$90 \$511 \$3 NWELL \$502 PWELL CLKBUF_X1
X$91 \$3 NWELL PWELL FILLCELL_X1
X$92 \$494 \$3 NWELL PWELL LOGIC0_X1
X$93 \$3 NWELL PWELL FILLCELL_X8
X$94 \$3 NWELL PWELL FILLCELL_X2
X$95 \$746 \$3 NWELL \$552 PWELL CLKBUF_X1
X$96 \$3 NWELL PWELL FILLCELL_X2
X$97 \$197 \$554 \$176 NWELL \$732 \$3 PWELL OAI21_X1
X$98 \$3 NWELL PWELL FILLCELL_X2
X$99 \$554 \$222 NWELL \$746 \$3 PWELL XOR2_X2
X$100 \$427 \$3 NWELL \$479 PWELL CLKBUF_X1
X$101 \$197 \$554 NWELL \$3 \$238 PWELL XNOR2_X1
X$102 \$3 NWELL PWELL FILLCELL_X4
X$103 \$430 \$428 \$502 \$429 \$63 NWELL \$3 \$555 PWELL OAI221_X1
X$104 \$3 NWELL PWELL FILLCELL_X4
X$105 \$3 NWELL PWELL FILLCELL_X2
X$106 \$371 \$197 \$554 \$3 \$750 NWELL PWELL AOI21_X1
X$107 \$3 NWELL PWELL FILLCELL_X1
X$108 \$245 \$3 NWELL \$781 PWELL CLKBUF_X1
X$109 \$3 NWELL PWELL NWELL TAPCELL_X1
X$110 \$3 NWELL PWELL FILLCELL_X1
X$111 \$753 \$3 NWELL \$482 PWELL CLKBUF_X1
X$112 \$626 \$482 \$758 \$557 NWELL \$3 \$744 PWELL OAI22_X1
X$113 \$737 \$557 \$479 \$3 NWELL \$741 PWELL MUX2_X1
X$114 \$494 \$557 \$482 \$3 NWELL \$490 PWELL MUX2_X1
X$115 \$3 NWELL PWELL FILLCELL_X1
X$116 \$3 NWELL PWELL FILLCELL_X2
X$117 NWELL VIA_via1_2_940_340_1_3_300_300
X$118 NWELL VIA_via2_3_940_340_1_3_320_320
X$119 NWELL VIA_via3_4_940_340_1_3_320_320
X$120 \$3 \$735 \$431 \$720 NWELL PWELL DFF_X2
X$121 \$3 NWELL PWELL FILLCELL_X8
X$122 \$3 \$627 \$431 \$573 NWELL PWELL DFF_X2
X$123 \$3 NWELL PWELL FILLCELL_X2
X$124 \$3 NWELL PWELL FILLCELL_X16
X$125 \$487 \$3 NWELL \$486 PWELL CLKBUF_X1
X$126 \$3 NWELL PWELL FILLCELL_X1
X$127 \$3 NWELL PWELL FILLCELL_X8
X$128 \$3 NWELL PWELL FILLCELL_X4
X$129 \$486 \$3 NWELL \$572 PWELL CLKBUF_X1
X$130 \$3 NWELL PWELL FILLCELL_X8
X$131 \$3 NWELL PWELL NWELL TAPCELL_X1
X$132 \$3 NWELL PWELL FILLCELL_X16
X$133 \$3 NWELL PWELL FILLCELL_X4
X$134 \$558 \$3 NWELL \$559 PWELL CLKBUF_X1
X$135 \$3 NWELL PWELL FILLCELL_X2
X$136 \$3 NWELL PWELL FILLCELL_X2
X$137 \$3 NWELL PWELL FILLCELL_X1
X$138 \$573 \$3 NWELL \$710 PWELL CLKBUF_X1
X$139 \$3 NWELL PWELL FILLCELL_X8
X$140 \$3 NWELL PWELL FILLCELL_X4
X$141 NWELL VIA_via1_2_940_340_1_3_300_300
X$142 NWELL VIA_via2_3_940_340_1_3_320_320
X$143 NWELL VIA_via3_4_940_340_1_3_320_320
X$144 \$710 \$3 NWELL \$558 PWELL CLKBUF_X1
X$145 \$3 NWELL PWELL FILLCELL_X16
X$146 \$3 NWELL PWELL FILLCELL_X1
X$147 \$691 \$3 NWELL zero_flag PWELL CLKBUF_X1
X$148 \$572 \$3 NWELL \$680 PWELL CLKBUF_X1
X$149 \$686 \$3 NWELL \$691 PWELL CLKBUF_X1
X$150 \$3 NWELL PWELL FILLCELL_X2
X$151 \$680 \$3 NWELL result[7] PWELL CLKBUF_X1
X$152 \$3 NWELL PWELL NWELL TAPCELL_X1
X$153 \$3 NWELL PWELL NWELL TAPCELL_X1
X$154 \$162 \$1153 \$1111 NWELL \$1151 \$3 PWELL OAI21_X1
X$155 \$3 NWELL PWELL FILLCELL_X1
X$156 \$3 NWELL PWELL FILLCELL_X1
X$157 \$1151 \$3 NWELL \$1084 PWELL INV_X1
X$158 \$1042 \$3 NWELL \$839 PWELL CLKBUF_X1
X$159 \$775 \$1112 \$1084 \$1004 \$1055 NWELL \$3 PWELL AOI211_X2
X$160 \$1142 \$1002 \$1111 \$3 \$1078 NWELL PWELL AOI21_X1
X$161 \$3 NWELL PWELL FILLCELL_X2
X$162 \$1101 \$366 \$1185 \$1208 NWELL \$1184 \$3 PWELL OAI211_X1
X$163 \$176 \$1137 \$3 NWELL \$1208 PWELL NAND2_X1
X$164 \$1184 \$3 NWELL \$1112 PWELL CLKBUF_X1
X$165 \$3 NWELL PWELL FILLCELL_X16
X$166 \$3 NWELL PWELL FILLCELL_X2
X$167 rst_n \$3 NWELL \$869 PWELL CLKBUF_X2
X$168 \$3 NWELL PWELL FILLCELL_X4
X$169 \$3 NWELL PWELL FILLCELL_X1
X$170 \$1113 \$839 NWELL \$3 \$1186 PWELL AND2_X1
X$171 \$3 NWELL PWELL FILLCELL_X1
X$172 \$1055 \$3 NWELL \$1006 PWELL CLKBUF_X1
X$173 \$1078 \$3 NWELL \$1115 PWELL CLKBUF_X1
X$174 \$1056 \$3 NWELL \$1114 PWELL CLKBUF_X1
X$175 \$921 \$3 NWELL \$1113 PWELL INV_X1
X$176 \$869 \$3 NWELL \$557 PWELL BUF_X2
X$177 \$921 \$557 \$1115 \$3 \$1059 NWELL PWELL AOI21_X1
X$178 \$3 \$1123 \$1116 \$1121 NWELL PWELL DFF_X2
X$179 \$1070 \$3 NWELL \$1123 PWELL CLKBUF_X1
X$180 \$3 NWELL PWELL FILLCELL_X8
X$181 \$3 NWELL PWELL FILLCELL_X4
X$182 \$1121 \$3 NWELL \$1067 PWELL CLKBUF_X1
X$183 \$3 NWELL PWELL FILLCELL_X4
X$184 \$3 NWELL PWELL FILLCELL_X2
X$185 \$3 NWELL PWELL FILLCELL_X2
X$186 \$3 NWELL PWELL NWELL TAPCELL_X1
X$187 \$1113 \$1114 NWELL \$3 \$1319 PWELL AND2_X1
X$188 \$3 NWELL PWELL FILLCELL_X2
X$189 \$3 \$1187 \$1116 \$1195 NWELL PWELL DFF_X2
X$190 \$3 NWELL PWELL FILLCELL_X16
X$191 \$1195 \$3 NWELL \$1188 PWELL CLKBUF_X1
X$192 \$3 NWELL PWELL FILLCELL_X4
X$193 \$3 NWELL PWELL FILLCELL_X2
X$194 \$1193 \$3 NWELL \$1062 PWELL CLKBUF_X1
X$195 \$1265 \$3 NWELL \$1061 PWELL CLKBUF_X1
X$196 \$1188 \$3 NWELL \$855 PWELL CLKBUF_X1
X$197 \$3 NWELL PWELL FILLCELL_X1
X$198 \$3 NWELL PWELL FILLCELL_X16
X$199 \$3 NWELL PWELL FILLCELL_X1
X$200 \$3 NWELL PWELL NWELL TAPCELL_X1
X$201 \$3 NWELL PWELL FILLCELL_X16
X$202 \$3 NWELL PWELL FILLCELL_X8
X$203 \$3 NWELL PWELL FILLCELL_X1
X$204 \$3 NWELL PWELL NWELL TAPCELL_X1
X$205 \$3 NWELL PWELL FILLCELL_X32
X$206 \$3 NWELL PWELL FILLCELL_X8
X$207 \$3 NWELL PWELL FILLCELL_X4
X$208 \$3 NWELL PWELL FILLCELL_X2
X$209 \$3 NWELL PWELL FILLCELL_X1
X$210 \$3 NWELL PWELL NWELL TAPCELL_X1
X$211 NWELL VIA_via1_2_940_340_1_3_300_300
X$212 NWELL VIA_via2_3_940_340_1_3_320_320
X$213 NWELL VIA_via3_4_940_340_1_3_320_320
X$214 NWELL VIA_via1_2_940_340_1_3_300_300
X$215 NWELL VIA_via2_3_940_340_1_3_320_320
X$216 NWELL VIA_via3_4_940_340_1_3_320_320
X$217 NWELL VIA_via1_2_940_340_1_3_300_300
X$218 NWELL VIA_via2_3_940_340_1_3_320_320
X$219 NWELL VIA_via3_4_940_340_1_3_320_320
X$220 \$720 \$3 NWELL \$714 PWELL CLKBUF_X1
X$221 \$3 NWELL PWELL FILLCELL_X1
X$222 \$3 NWELL PWELL FILLCELL_X8
X$223 \$3 NWELL PWELL FILLCELL_X4
X$224 \$714 \$3 NWELL \$686 PWELL CLKBUF_X1
X$225 \$3 NWELL PWELL FILLCELL_X8
X$226 \$3 NWELL PWELL FILLCELL_X1
X$227 \$3 NWELL PWELL NWELL TAPCELL_X1
X$228 \$3 NWELL PWELL FILLCELL_X8
X$229 \$3 NWELL PWELL FILLCELL_X2
X$230 \$3 NWELL PWELL FILLCELL_X8
X$231 \$741 \$3 NWELL \$627 PWELL CLKBUF_X1
X$232 \$3 NWELL PWELL FILLCELL_X2
X$233 \$3 NWELL PWELL FILLCELL_X1
X$234 \$3 \$844 \$431 \$857 NWELL PWELL DFF_X2
X$235 \$3 NWELL PWELL FILLCELL_X8
X$236 \$803 \$3 NWELL \$431 PWELL CLKBUF_X3
X$237 \$3 NWELL PWELL FILLCELL_X2
X$238 \$3 NWELL PWELL FILLCELL_X16
X$239 \$3 NWELL PWELL FILLCELL_X8
X$240 \$3 NWELL PWELL FILLCELL_X4
X$241 NWELL VIA_via1_2_940_340_1_3_300_300
X$242 NWELL VIA_via2_3_940_340_1_3_320_320
X$243 NWELL VIA_via3_4_940_340_1_3_320_320
X$244 \$856 \$3 NWELL \$795 PWELL CLKBUF_X1
X$245 \$3 NWELL PWELL FILLCELL_X16
X$246 \$849 \$3 NWELL result[5] PWELL CLKBUF_X1
X$247 \$689 \$3 NWELL result[3] PWELL CLKBUF_X1
X$248 \$559 \$3 NWELL result[4] PWELL CLKBUF_X1
X$249 \$629 \$3 NWELL result[0] PWELL CLKBUF_X1
X$250 \$795 \$3 NWELL \$689 PWELL CLKBUF_X1
X$251 \$630 \$3 NWELL result[1] PWELL CLKBUF_X1
X$252 \$3 NWELL PWELL NWELL TAPCELL_X1
X$253 \$926 \$3 NWELL overflow_flag PWELL CLKBUF_X1
X$254 \$850 \$3 NWELL result[6] PWELL CLKBUF_X1
X$255 \$845 \$3 NWELL result[2] PWELL CLKBUF_X1
X$256 \$783 \$3 NWELL \$849 PWELL CLKBUF_X1
X$257 \$3 NWELL PWELL NWELL TAPCELL_X1
X$258 \$1162 \$3 NWELL \$996 PWELL INV_X1
X$259 \$1162 \$893 \$3 NWELL \$1222 PWELL NAND2_X1
X$260 \$3 NWELL PWELL FILLCELL_X1
X$261 \$896 a[1] NWELL \$1097 \$3 PWELL XOR2_X2
X$262 \$3 NWELL PWELL FILLCELL_X1
X$263 \$1097 \$224 \$996 \$3 \$1182 NWELL PWELL AOI21_X2
X$264 \$1217 \$1270 \$1076 \$1230 \$1279 \$3 NWELL \$1171 PWELL AOI221_X1
X$265 \$3 NWELL PWELL FILLCELL_X4
X$266 \$3 NWELL PWELL FILLCELL_X1
X$267 \$1097 \$233 \$1220 \$335 \$1096 \$3 NWELL \$1225 PWELL AOI221_X1
X$268 \$3 NWELL PWELL FILLCELL_X2
X$269 \$3 NWELL PWELL FILLCELL_X16
X$270 \$3 NWELL PWELL NWELL TAPCELL_X1
X$271 \$3 NWELL PWELL FILLCELL_X4
X$272 \$3 NWELL PWELL FILLCELL_X2
X$273 \$3 NWELL PWELL NWELL TAPCELL_X1
X$274 \$3 NWELL PWELL FILLCELL_X32
X$275 NWELL VIA_via1_2_940_340_1_3_300_300
X$276 NWELL VIA_via2_3_940_340_1_3_320_320
X$277 NWELL VIA_via3_4_940_340_1_3_320_320
X$278 \$3 NWELL PWELL FILLCELL_X4
X$279 \$3 NWELL PWELL FILLCELL_X2
X$280 \$3 NWELL PWELL FILLCELL_X1
X$281 \$1097 \$1222 NWELL \$3 \$1270 PWELL XNOR2_X1
X$282 \$1097 \$996 \$893 \$3 NWELL \$1279 PWELL NAND3_X1
X$283 \$3 NWELL PWELL FILLCELL_X8
X$284 \$3 NWELL PWELL FILLCELL_X4
X$285 \$3 NWELL PWELL FILLCELL_X2
X$286 \$3 NWELL PWELL FILLCELL_X1
X$287 \$3 NWELL PWELL NWELL TAPCELL_X1
X$288 \$1254 \$825 \$1253 \$3 \$356 NWELL PWELL NAND3_X4
X$289 opcode[1] \$1254 \$3 NWELL \$227 PWELL NAND2_X2
X$290 opcode[1] \$1261 \$3 NWELL \$999 PWELL NAND2_X2
X$291 \$913 \$1108 \$1261 \$1258 NWELL \$1178 \$3 PWELL OAI211_X1
X$292 \$913 \$1182 \$1177 \$3 NWELL \$1246 PWELL OR3_X1
X$293 \$1246 \$1258 \$919 \$1254 \$3 NWELL \$1242 PWELL NAND4_X1
X$294 \$1258 \$1254 \$3 NWELL \$63 PWELL NAND2_X2
X$295 \$63 \$1182 \$3 NWELL \$1230 PWELL NOR2_X1
X$296 \$233 \$1258 \$1101 \$1137 NWELL \$1298 \$3 PWELL OAI211_X1
X$297 \$1258 \$1261 \$3 NWELL \$294 PWELL NAND2_X2
X$298 \$1298 \$3 NWELL \$1185 PWELL CLKBUF_X1
X$299 \$3 NWELL PWELL FILLCELL_X16
X$300 \$3 NWELL PWELL FILLCELL_X8
X$301 \$3 NWELL PWELL FILLCELL_X2
X$302 \$123 opcode[1] \$1305 \$3 NWELL \$1217 PWELL NOR3_X1
X$303 NWELL VIA_via1_2_940_340_1_3_300_300
X$304 NWELL VIA_via2_3_940_340_1_3_320_320
X$305 NWELL VIA_via3_4_940_340_1_3_320_320
X$306 \$998 opcode[1] \$3 NWELL \$1253 PWELL NOR2_X2
X$307 \$3 NWELL PWELL FILLCELL_X2
X$308 \$3 \$1254 opcode[1] \$1050 \$233 NWELL PWELL NOR3_X4
X$309 \$123 opcode[1] \$3 NWELL \$1258 PWELL NOR2_X2
X$310 \$3 NWELL PWELL FILLCELL_X8
X$311 \$1254 \$3 NWELL \$1261 PWELL INV_X1
X$312 \$3 NWELL PWELL FILLCELL_X32
X$313 NWELL VIA_via1_2_940_340_1_3_300_300
X$314 NWELL VIA_via2_3_940_340_1_3_320_320
X$315 NWELL VIA_via3_4_940_340_1_3_320_320
X$316 \$3 NWELL PWELL FILLCELL_X16
X$317 \$3 \$1291 \$1116 \$1283 NWELL PWELL DFF_X2
X$318 \$1186 \$3 NWELL \$1291 PWELL CLKBUF_X1
X$319 \$1059 \$3 NWELL \$1187 PWELL CLKBUF_X1
X$320 \$3 NWELL PWELL FILLCELL_X8
X$321 \$3 NWELL PWELL FILLCELL_X4
X$322 \$3 NWELL PWELL FILLCELL_X2
X$323 \$3 NWELL PWELL FILLCELL_X4
X$324 \$3 NWELL PWELL NWELL TAPCELL_X1
X$325 \$3 \$1320 \$1116 \$1339 NWELL PWELL DFF_X2
X$326 NWELL VIA_via1_2_940_340_1_3_300_300
X$327 NWELL VIA_via2_3_940_340_1_3_320_320
X$328 NWELL VIA_via3_4_940_340_1_3_320_320
X$329 \$803 \$3 NWELL \$1116 PWELL CLKBUF_X3
X$330 \$3 NWELL PWELL FILLCELL_X8
X$331 \$3 NWELL PWELL FILLCELL_X32
X$332 \$1283 \$3 NWELL \$1193 PWELL CLKBUF_X1
X$333 \$3 NWELL PWELL FILLCELL_X8
X$334 \$3 NWELL PWELL FILLCELL_X2
X$335 \$3 NWELL PWELL FILLCELL_X4
X$336 \$1339 \$3 NWELL \$1265 PWELL CLKBUF_X1
X$337 \$3 NWELL PWELL FILLCELL_X32
X$338 NWELL VIA_via1_2_940_340_1_3_300_300
X$339 NWELL VIA_via2_3_940_340_1_3_320_320
X$340 NWELL VIA_via3_4_940_340_1_3_320_320
X$341 \$3 NWELL PWELL FILLCELL_X32
X$342 \$3 NWELL PWELL FILLCELL_X16
X$343 \$3 NWELL PWELL NWELL TAPCELL_X1
X$344 \$3 NWELL PWELL FILLCELL_X8
X$345 \$3 NWELL PWELL FILLCELL_X1
X$346 \$3 NWELL PWELL NWELL TAPCELL_X1
X$347 \$3 NWELL PWELL NWELL TAPCELL_X1
X$348 NWELL VIA_via5_6_940_960_2_2_600_600
X$349 NWELL VIA_via4_5_940_960_2_2_600_600
X$350 NWELL VIA_via6_7_940_960_1_1_600_600
X$351 NWELL VIA_via5_6_940_960_2_2_600_600
X$352 NWELL VIA_via4_5_940_960_2_2_600_600
X$353 NWELL VIA_via6_7_940_960_1_1_600_600
X$354 NWELL VIA_via5_6_940_960_2_2_600_600
X$355 NWELL VIA_via4_5_940_960_2_2_600_600
X$356 NWELL VIA_via6_7_940_960_1_1_600_600
X$357 NWELL VIA_via5_6_940_960_2_2_600_600
X$358 NWELL VIA_via4_5_940_960_2_2_600_600
X$359 NWELL VIA_via6_7_940_960_1_1_600_600
X$360 NWELL VIA_via5_6_940_960_2_2_600_600
X$361 NWELL VIA_via4_5_940_960_2_2_600_600
X$362 NWELL VIA_via6_7_940_960_1_1_600_600
X$363 NWELL VIA_via5_6_940_960_2_2_600_600
X$364 NWELL VIA_via4_5_940_960_2_2_600_600
X$365 NWELL VIA_via6_7_940_960_1_1_600_600
X$366 NWELL VIA_via5_6_940_960_2_2_600_600
X$367 NWELL VIA_via4_5_940_960_2_2_600_600
X$368 NWELL VIA_via6_7_940_960_1_1_600_600
X$369 NWELL VIA_via5_6_940_960_2_2_600_600
X$370 NWELL VIA_via4_5_940_960_2_2_600_600
X$371 NWELL VIA_via6_7_940_960_1_1_600_600
X$372 NWELL VIA_via5_6_940_960_2_2_600_600
X$373 NWELL VIA_via4_5_940_960_2_2_600_600
X$374 NWELL VIA_via6_7_940_960_1_1_600_600
X$375 NWELL VIA_via5_6_940_960_2_2_600_600
X$376 NWELL VIA_via4_5_940_960_2_2_600_600
X$377 NWELL VIA_via6_7_940_960_1_1_600_600
X$378 NWELL VIA_via5_6_940_960_2_2_600_600
X$379 NWELL VIA_via4_5_940_960_2_2_600_600
X$380 NWELL VIA_via6_7_940_960_1_1_600_600
X$381 NWELL VIA_via5_6_940_960_2_2_600_600
X$382 NWELL VIA_via4_5_940_960_2_2_600_600
X$383 NWELL VIA_via6_7_940_960_1_1_600_600
X$384 NWELL VIA_via5_6_940_960_2_2_600_600
X$385 NWELL VIA_via4_5_940_960_2_2_600_600
X$386 NWELL VIA_via6_7_940_960_1_1_600_600
X$387 NWELL VIA_via5_6_940_960_2_2_600_600
X$388 NWELL VIA_via4_5_940_960_2_2_600_600
X$389 NWELL VIA_via6_7_940_960_1_1_600_600
X$390 NWELL VIA_via5_6_940_960_2_2_600_600
X$391 NWELL VIA_via4_5_940_960_2_2_600_600
X$392 NWELL VIA_via6_7_940_960_1_1_600_600
X$393 NWELL VIA_via5_6_940_960_2_2_600_600
X$394 NWELL VIA_via4_5_940_960_2_2_600_600
X$395 NWELL VIA_via6_7_940_960_1_1_600_600
X$396 NWELL VIA_via5_6_940_960_2_2_600_600
X$397 NWELL VIA_via4_5_940_960_2_2_600_600
X$398 NWELL VIA_via6_7_940_960_1_1_600_600
X$399 NWELL VIA_via5_6_940_960_2_2_600_600
X$400 NWELL VIA_via4_5_940_960_2_2_600_600
X$401 NWELL VIA_via6_7_940_960_1_1_600_600
X$402 NWELL VIA_via5_6_940_960_2_2_600_600
X$403 NWELL VIA_via4_5_940_960_2_2_600_600
X$404 NWELL VIA_via6_7_940_960_1_1_600_600
X$405 NWELL VIA_via5_6_940_960_2_2_600_600
X$406 NWELL VIA_via4_5_940_960_2_2_600_600
X$407 NWELL VIA_via6_7_940_960_1_1_600_600
X$408 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$409 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$410 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$411 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$412 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$413 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$414 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$415 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$416 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$417 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$418 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$419 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$420 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$421 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$422 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$423 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$424 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$425 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$426 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$427 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$428 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$429 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$430 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$431 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$432 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$433 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$434 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$435 NWELL VIA_via9_10_1600_2400_1_1_3360_3360
X$436 NWELL VIA_via8_9_1600_1600_1_1_1680_1680
X$437 NWELL VIA_via7_8_1600_960_1_1_1680_1680
X$438 \$3 NWELL PWELL FILLCELL_X16
X$439 \$3 NWELL PWELL NWELL TAPCELL_X1
X$440 \$3 NWELL PWELL FILLCELL_X2
X$441 \$3 NWELL PWELL NWELL TAPCELL_X1
X$442 \$3 NWELL PWELL FILLCELL_X8
X$443 \$3 NWELL PWELL FILLCELL_X4
X$444 \$991 a[2] \$893 \$3 \$993 NWELL PWELL AOI21_X1
X$445 NWELL VIA_via1_2_940_340_1_3_300_300
X$446 NWELL VIA_via2_3_940_340_1_3_320_320
X$447 NWELL VIA_via3_4_940_340_1_3_320_320
X$448 \$931 \$279 \$993 \$3 \$1076 NWELL PWELL AOI21_X1
X$449 \$279 \$351 \$827 NWELL \$931 \$3 PWELL OAI21_X1
X$450 \$3 NWELL PWELL FILLCELL_X1
X$451 \$3 NWELL PWELL FILLCELL_X2
X$452 \$3 NWELL PWELL FILLCELL_X4
X$453 \$3 NWELL PWELL FILLCELL_X1
X$454 \$996 \$893 \$3 NWELL \$895 PWELL NOR2_X1
X$455 \$893 a[1] \$895 \$896 \$3 \$858 NWELL PWELL AOI211_X1
X$456 \$3 NWELL PWELL FILLCELL_X1
X$457 \$3 NWELL PWELL FILLCELL_X1
X$458 \$896 \$574 \$357 \$858 \$3 \$861 NWELL PWELL AOI211_X1
X$459 \$284 \$3 NWELL \$1019 PWELL BUF_X2
X$460 \$895 \$896 \$3 NWELL \$801 PWELL NAND2_X1
X$461 \$3 NWELL PWELL FILLCELL_X1
X$462 \$811 \$255 NWELL \$3 \$903 PWELL AND2_X1
X$463 \$861 \$819 \$903 \$3 NWELL \$775 PWELL OR3_X1
X$464 \$606 \$356 \$769 \$3 NWELL \$904 PWELL NOR3_X1
X$465 \$284 \$3 NWELL \$769 PWELL BUF_X1
X$466 \$3 NWELL PWELL FILLCELL_X4
X$467 \$3 NWELL PWELL FILLCELL_X2
X$468 \$3 NWELL PWELL FILLCELL_X4
X$469 \$3 NWELL PWELL FILLCELL_X1
X$470 \$1019 NWELL \$896 \$3 PWELL BUF_X4
X$471 \$996 \$896 \$893 \$3 NWELL \$811 PWELL NOR3_X1
X$472 \$3 NWELL PWELL FILLCELL_X8
X$473 \$3 NWELL PWELL FILLCELL_X1
X$474 \$904 \$1077 \$287 \$3 \$1098 NWELL PWELL AOI21_X1
X$475 \$3 NWELL PWELL FILLCELL_X4
X$476 \$825 \$998 \$999 \$3 NWELL \$770 PWELL OR3_X1
X$477 NWELL VIA_via1_2_940_340_1_3_300_300
X$478 NWELL VIA_via2_3_940_340_1_3_320_320
X$479 NWELL VIA_via3_4_940_340_1_3_320_320
X$480 b[2] \$998 \$999 \$3 NWELL \$357 PWELL OR3_X2
X$481 \$772 \$818 \$3 NWELL \$255 PWELL NOR2_X2
X$482 \$3 NWELL PWELL FILLCELL_X1
X$483 \$3 NWELL PWELL FILLCELL_X1
X$484 \$825 a[2] \$3 NWELL \$918 PWELL NAND2_X1
X$485 \$3 NWELL PWELL NWELL TAPCELL_X1
X$486 \$3 NWELL PWELL FILLCELL_X2
X$487 \$3 \$818 \$1050 \$999 \$827 NWELL PWELL NOR3_X4
X$488 \$909 \$366 \$869 \$960 NWELL \$972 \$3 PWELL OAI211_X1
X$489 b[2] a[2] \$3 NWELL \$909 PWELL NAND2_X1
X$490 \$794 \$827 \$972 \$233 \$833 \$973 NWELL \$3 PWELL AOI221_X2
X$491 \$914 \$909 NWELL \$3 \$833 PWELL AND2_X1
X$492 \$3 NWELL PWELL FILLCELL_X2
X$493 \$3 NWELL PWELL FILLCELL_X1
X$494 \$255 \$230 \$1089 \$1088 \$176 \$3 NWELL \$1046 PWELL AOI221_X1
X$495 \$3 NWELL PWELL FILLCELL_X4
X$496 \$3 NWELL PWELL FILLCELL_X1
X$497 \$909 \$914 \$3 NWELL \$913 PWELL NAND2_X2
X$498 \$973 \$1046 \$1109 \$3 NWELL \$1042 PWELL NAND3_X1
X$499 \$549 \$918 \$919 NWELL \$3 \$777 PWELL AND3_X1
X$500 \$3 NWELL PWELL FILLCELL_X1
X$501 \$3 \$62 \$549 \$919 \$918 NWELL PWELL AOI21_X4
X$502 \$3 NWELL PWELL FILLCELL_X4
X$503 \$3 NWELL PWELL FILLCELL_X1
X$504 \$957 \$3 NWELL PWELL LOGIC0_X1
X$505 \$3 NWELL PWELL FILLCELL_X16
X$506 \$750 \$3 NWELL \$975 PWELL CLKBUF_X1
X$507 \$980 \$3 NWELL \$780 PWELL CLKBUF_X1
X$508 \$3 NWELL PWELL FILLCELL_X2
X$509 \$895 \$549 \$3 NWELL \$1001 PWELL NOR2_X1
X$510 \$3 NWELL PWELL FILLCELL_X16
X$511 NWELL VIA_via1_2_940_340_1_3_300_300
X$512 NWELL VIA_via2_3_940_340_1_3_320_320
X$513 NWELL VIA_via3_4_940_340_1_3_320_320
X$514 \$3 NWELL PWELL FILLCELL_X8
X$515 \$3 NWELL PWELL FILLCELL_X2
X$516 \$3 NWELL PWELL FILLCELL_X1
X$517 \$1003 \$295 NWELL \$3 \$1002 PWELL AND2_X1
X$518 \$63 \$1004 \$869 \$975 \$294 NWELL \$3 \$1056 PWELL OAI221_X1
X$519 \$295 \$1003 \$3 NWELL \$1004 PWELL NAND2_X1
X$520 \$3 NWELL PWELL FILLCELL_X4
X$521 \$3 NWELL PWELL FILLCELL_X2
X$522 \$3 NWELL PWELL FILLCELL_X1
X$523 \$866 \$781 \$1115 \$1006 \$3 NWELL \$626 PWELL NAND4_X1
X$524 \$869 \$840 \$3 NWELL \$921 PWELL NOR2_X2
X$525 \$921 \$557 \$781 \$3 \$841 NWELL PWELL AOI21_X1
X$526 \$921 \$557 \$860 \$3 \$842 NWELL PWELL AOI21_X1
X$527 \$3 NWELL PWELL FILLCELL_X2
X$528 \$3 NWELL PWELL NWELL TAPCELL_X1
X$529 \$3 NWELL PWELL FILLCELL_X4
X$530 \$3 NWELL PWELL FILLCELL_X2
X$531 \$3 NWELL PWELL FILLCELL_X1
X$532 \$921 \$557 \$1006 \$3 \$1070 NWELL PWELL AOI21_X1
X$533 \$3 NWELL PWELL FILLCELL_X2
X$534 \$841 \$3 NWELL \$1016 PWELL CLKBUF_X1
X$535 NWELL VIA_via1_2_940_340_1_3_300_300
X$536 NWELL VIA_via2_3_940_340_1_3_320_320
X$537 NWELL VIA_via3_4_940_340_1_3_320_320
X$538 clk \$3 NWELL \$803 PWELL CLKBUF_X3
X$539 \$842 \$3 NWELL \$948 PWELL CLKBUF_X1
X$540 \$843 \$3 NWELL \$844 PWELL CLKBUF_X1
X$541 \$3 \$948 \$431 \$946 NWELL PWELL DFF_X2
X$542 \$3 NWELL PWELL FILLCELL_X8
X$543 \$3 NWELL PWELL FILLCELL_X4
X$544 \$3 NWELL PWELL FILLCELL_X1
X$545 \$946 \$3 NWELL \$939 PWELL CLKBUF_X1
X$546 \$857 \$3 NWELL \$856 PWELL CLKBUF_X1
X$547 \$3 NWELL PWELL FILLCELL_X8
X$548 \$3 NWELL PWELL FILLCELL_X1
X$549 \$939 \$3 NWELL \$783 PWELL CLKBUF_X1
X$550 \$3 NWELL PWELL FILLCELL_X2
X$551 \$3 \$1016 \$431 \$1015 NWELL PWELL DFF_X2
X$552 \$3 NWELL PWELL FILLCELL_X8
X$553 \$3 NWELL PWELL FILLCELL_X4
X$554 \$3 NWELL PWELL FILLCELL_X2
X$555 \$1015 \$3 NWELL \$1012 PWELL CLKBUF_X1
X$556 \$3 NWELL PWELL FILLCELL_X4
X$557 \$3 NWELL PWELL FILLCELL_X2
X$558 \$1067 \$3 NWELL \$925 PWELL CLKBUF_X1
X$559 \$3 NWELL PWELL FILLCELL_X2
X$560 NWELL VIA_via1_2_940_340_1_3_300_300
X$561 NWELL VIA_via2_3_940_340_1_3_320_320
X$562 NWELL VIA_via3_4_940_340_1_3_320_320
X$563 \$3 NWELL PWELL FILLCELL_X1
X$564 \$1012 \$3 NWELL \$1008 PWELL CLKBUF_X1
X$565 \$3 NWELL PWELL FILLCELL_X8
X$566 \$3 NWELL PWELL FILLCELL_X8
X$567 \$3 NWELL PWELL NWELL TAPCELL_X1
X$568 \$3 NWELL PWELL FILLCELL_X4
X$569 \$855 \$3 NWELL \$630 PWELL CLKBUF_X1
X$570 \$3 NWELL PWELL FILLCELL_X1
X$571 \$925 \$3 NWELL \$629 PWELL CLKBUF_X1
X$572 \$3 NWELL PWELL FILLCELL_X1
X$573 \$1008 \$3 NWELL \$850 PWELL CLKBUF_X1
X$574 \$3 NWELL PWELL FILLCELL_X2
X$575 \$3 NWELL PWELL FILLCELL_X4
X$576 \$3 NWELL PWELL FILLCELL_X1
X$577 \$1062 \$3 NWELL \$845 PWELL CLKBUF_X1
X$578 \$1061 \$3 NWELL \$926 PWELL CLKBUF_X1
X$579 \$3 NWELL PWELL FILLCELL_X8
X$580 \$3 NWELL PWELL FILLCELL_X4
X$581 \$3 NWELL PWELL NWELL TAPCELL_X1
X$582 \$3 NWELL PWELL NWELL TAPCELL_X1
X$583 \$3 NWELL PWELL FILLCELL_X8
X$584 \$3 NWELL PWELL NWELL TAPCELL_X1
X$585 \$3 NWELL PWELL FILLCELL_X4
X$586 \$3 NWELL PWELL FILLCELL_X2
X$587 \$3 NWELL PWELL NWELL TAPCELL_X1
X$588 \$3 NWELL PWELL FILLCELL_X2
X$589 \$3 NWELL PWELL FILLCELL_X1
X$590 b[6] \$3 NWELL \$101 PWELL CLKBUF_X1
X$591 \$90 \$3 NWELL \$200 PWELL INV_X2
X$592 \$352 \$200 \$3 NWELL \$382 PWELL NOR2_X1
X$593 \$397 \$90 \$18 \$3 NWELL \$351 PWELL MUX2_X1
X$594 \$382 \$200 \$18 \$3 \$215 NWELL PWELL AOI21_X1
X$595 a[6] \$3 NWELL \$131 PWELL CLKBUF_X1
X$596 \$3 NWELL PWELL FILLCELL_X1
X$597 \$279 \$215 NWELL \$3 \$280 PWELL AND2_X1
X$598 \$217 \$3 NWELL \$305 PWELL BUF_X1
X$599 a[4] \$3 NWELL \$217 PWELL CLKBUF_X1
X$600 \$3 NWELL PWELL FILLCELL_X4
X$601 \$3 NWELL PWELL FILLCELL_X2
X$602 \$305 NWELL \$18 \$3 PWELL BUF_X4
X$603 \$280 \$356 \$173 \$354 \$326 NWELL \$3 PWELL AOI211_X2
X$604 \$278 \$356 \$279 \$306 \$394 NWELL \$3 PWELL AOI211_X2
X$605 \$3 NWELL PWELL FILLCELL_X1
X$606 \$173 \$306 \$172 \$356 \$3 \$220 NWELL PWELL AOI211_X1
X$607 \$3 NWELL PWELL FILLCELL_X1
X$608 \$128 \$284 \$149 NWELL \$3 \$287 PWELL OAI21_X2
X$609 \$3 NWELL PWELL FILLCELL_X1
X$610 \$222 \$3 NWELL \$325 PWELL BUF_X2
X$611 \$3 NWELL PWELL FILLCELL_X1
X$612 \$129 \$67 \$197 \$3 \$289 NWELL PWELL AOI21_X2
X$613 \$224 \$3 NWELL \$342 PWELL BUF_X1
X$614 \$3 NWELL PWELL FILLCELL_X8
X$615 \$3 NWELL PWELL FILLCELL_X1
X$616 \$3 NWELL PWELL NWELL TAPCELL_X1
X$617 \$233 \$26 \$225 \$335 \$56 \$339 NWELL \$3 PWELL AOI221_X2
X$618 \$231 \$230 \$396 \$176 \$134 \$265 NWELL \$3 PWELL AOI221_X2
X$619 \$321 \$104 \$233 \$3 \$203 NWELL PWELL AOI21_X1
X$620 \$3 NWELL PWELL FILLCELL_X2
X$621 \$357 \$173 \$149 \$3 \$416 NWELL PWELL AOI21_X1
X$622 \$3 NWELL PWELL FILLCELL_X2
X$623 \$3 NWELL PWELL FILLCELL_X1
X$624 \$325 NWELL \$197 \$3 PWELL BUF_X4
X$625 \$394 \$359 \$287 \$360 \$324 NWELL \$3 PWELL AOI211_X2
X$626 \$289 \$357 \$174 \$3 NWELL \$321 PWELL NOR3_X1
X$627 \$342 \$3 NWELL \$67 PWELL BUF_X2
X$628 \$599 \$339 \$3 NWELL \$359 PWELL NAND2_X1
X$629 \$3 NWELL PWELL FILLCELL_X4
X$630 \$3 NWELL PWELL FILLCELL_X2
X$631 \$3 NWELL PWELL FILLCELL_X1
X$632 \$366 \$103 \$3 NWELL \$396 PWELL NOR2_X1
X$633 \$397 b[3] NWELL \$3 \$458 PWELL AND2_X1
X$634 \$3 NWELL PWELL FILLCELL_X2
X$635 b[3] \$352 \$3 NWELL \$42 PWELL NOR2_X2
X$636 \$3 NWELL PWELL FILLCELL_X4
X$637 \$3 NWELL PWELL FILLCELL_X2
X$638 \$3 NWELL PWELL FILLCELL_X1
X$639 \$258 \$3 NWELL \$390 PWELL CLKBUF_X1
X$640 \$3 NWELL PWELL FILLCELL_X1
X$641 \$233 \$20 \$291 \$326 \$3 \$258 NWELL PWELL AOI211_X1
X$642 \$180 \$366 \$254 NWELL \$365 \$3 PWELL OAI21_X1
X$643 \$313 \$30 \$180 NWELL \$183 \$3 PWELL OAI21_X1
X$644 \$138 \$3 NWELL \$254 PWELL CLKBUF_X1
X$645 \$26 \$183 NWELL \$3 \$293 PWELL XNOR2_X1
X$646 \$3 NWELL PWELL FILLCELL_X16
X$647 \$238 \$103 \$240 NWELL \$3 \$430 PWELL AND3_X1
X$648 \$294 \$185 \$186 \$3 \$242 NWELL PWELL AOI21_X1
X$649 \$3 NWELL PWELL FILLCELL_X32
X$650 \$3 NWELL PWELL FILLCELL_X32
X$651 \$3 NWELL PWELL FILLCELL_X16
X$652 \$3 NWELL PWELL NWELL TAPCELL_X1
X$653 \$3 NWELL PWELL FILLCELL_X16
X$654 \$3 NWELL PWELL FILLCELL_X8
X$655 \$3 NWELL PWELL FILLCELL_X1
X$656 \$3 NWELL PWELL NWELL TAPCELL_X1
X$657 \$390 \$362 NWELL \$3 \$448 PWELL AND2_X1
X$658 \$30 \$313 NWELL \$3 \$292 PWELL XNOR2_X1
X$659 \$294 \$292 \$237 \$509 NWELL \$427 \$3 PWELL OAI211_X1
X$660 \$3 NWELL PWELL FILLCELL_X4
X$661 \$3 NWELL PWELL FILLCELL_X2
X$662 \$293 \$294 \$72 \$439 NWELL \$438 \$3 PWELL OAI211_X1
X$663 \$3 NWELL PWELL FILLCELL_X4
X$664 \$3 NWELL PWELL FILLCELL_X2
X$665 \$3 NWELL PWELL FILLCELL_X1
X$666 \$294 \$371 \$3 NWELL \$428 PWELL OR2_X1
X$667 \$552 \$374 NWELL \$3 \$429 PWELL XNOR2_X1
X$668 \$3 NWELL PWELL FILLCELL_X4
X$669 \$3 NWELL PWELL NWELL TAPCELL_X1
X$670 \$238 \$240 \$103 \$3 \$371 NWELL PWELL AOI21_X1
X$671 \$3 NWELL PWELL FILLCELL_X8
X$672 \$3 NWELL PWELL FILLCELL_X4
X$673 \$3 NWELL PWELL FILLCELL_X2
X$674 \$3 \$490 \$431 \$487 NWELL PWELL DFF_X2
X$675 \$3 NWELL PWELL FILLCELL_X32
X$676 \$3 NWELL PWELL FILLCELL_X32
X$677 \$3 NWELL PWELL FILLCELL_X2
X$678 \$3 NWELL PWELL NWELL TAPCELL_X1
X$679 NWELL VIA_via1_2_940_340_1_3_300_300
X$680 NWELL VIA_via5_6_940_960_2_2_600_600
X$681 NWELL VIA_via4_5_940_960_2_2_600_600
X$682 NWELL VIA_via6_7_940_960_1_1_600_600
X$683 NWELL VIA_via3_4_940_340_1_3_320_320
X$684 NWELL VIA_via2_3_940_340_1_3_320_320
X$685 NWELL VIA_via1_2_940_340_1_3_300_300
X$686 NWELL VIA_via5_6_940_960_2_2_600_600
X$687 NWELL VIA_via4_5_940_960_2_2_600_600
X$688 NWELL VIA_via6_7_940_960_1_1_600_600
X$689 NWELL VIA_via3_4_940_340_1_3_320_320
X$690 NWELL VIA_via2_3_940_340_1_3_320_320
X$691 NWELL VIA_via1_2_940_340_1_3_300_300
X$692 NWELL VIA_via5_6_940_960_2_2_600_600
X$693 NWELL VIA_via4_5_940_960_2_2_600_600
X$694 NWELL VIA_via6_7_940_960_1_1_600_600
X$695 NWELL VIA_via3_4_940_340_1_3_320_320
X$696 NWELL VIA_via2_3_940_340_1_3_320_320
X$697 NWELL VIA_via1_2_940_340_1_3_300_300
X$698 NWELL VIA_via5_6_940_960_2_2_600_600
X$699 NWELL VIA_via4_5_940_960_2_2_600_600
X$700 NWELL VIA_via6_7_940_960_1_1_600_600
X$701 NWELL VIA_via3_4_940_340_1_3_320_320
X$702 NWELL VIA_via2_3_940_340_1_3_320_320
X$703 NWELL VIA_via1_2_940_340_1_3_300_300
X$704 NWELL VIA_via5_6_940_960_2_2_600_600
X$705 NWELL VIA_via4_5_940_960_2_2_600_600
X$706 NWELL VIA_via6_7_940_960_1_1_600_600
X$707 NWELL VIA_via3_4_940_340_1_3_320_320
X$708 NWELL VIA_via2_3_940_340_1_3_320_320
X$709 \$3 NWELL PWELL FILLCELL_X8
X$710 \$3 NWELL PWELL NWELL TAPCELL_X1
X$711 \$3 NWELL PWELL FILLCELL_X4
X$712 \$3 NWELL PWELL FILLCELL_X2
X$713 \$3 NWELL PWELL NWELL TAPCELL_X1
X$714 \$3 NWELL PWELL FILLCELL_X16
X$715 \$3 NWELL PWELL FILLCELL_X1
X$716 \$224 \$3 NWELL \$893 PWELL BUF_X2
X$717 \$991 \$1127 \$3 NWELL \$606 PWELL NOR2_X1
X$718 \$893 \$1093 \$3 NWELL \$991 PWELL NOR2_X1
X$719 \$3 NWELL PWELL FILLCELL_X2
X$720 \$3 NWELL PWELL FILLCELL_X2
X$721 \$893 \$1162 NWELL \$3 \$1127 PWELL AND2_X1
X$722 a[1] \$3 NWELL \$1093 PWELL INV_X1
X$723 \$3 NWELL PWELL FILLCELL_X4
X$724 \$896 \$3 NWELL \$279 PWELL INV_X2
X$725 \$3 NWELL PWELL FILLCELL_X1
X$726 \$3 NWELL PWELL FILLCELL_X8
X$727 \$3 NWELL PWELL FILLCELL_X4
X$728 \$3 NWELL PWELL FILLCELL_X1
X$729 \$996 \$200 \$3 NWELL \$1137 PWELL NAND2_X1
X$730 \$3 NWELL PWELL FILLCELL_X16
X$731 \$999 \$1050 \$825 \$3 NWELL \$1077 PWELL NOR3_X1
X$732 \$3 NWELL PWELL FILLCELL_X4
X$733 b[2] \$3 NWELL \$825 PWELL INV_X2
X$734 \$3 NWELL PWELL FILLCELL_X2
X$735 \$3 NWELL PWELL FILLCELL_X2
X$736 \$3 NWELL PWELL FILLCELL_X1
X$737 a[1] \$896 NWELL \$3 \$1096 PWELL AND2_X1
X$738 \$3 NWELL PWELL FILLCELL_X2
X$739 \$3 NWELL PWELL FILLCELL_X1
X$740 \$1096 \$1127 \$1097 \$3 \$1108 NWELL PWELL AOI21_X2
X$741 \$896 \$1093 \$3 NWELL \$1177 PWELL NOR2_X1
X$742 \$279 \$1093 \$123 \$227 \$3 \$1220 NWELL PWELL AOI211_X1
X$743 \$1171 \$1098 \$1225 \$3 NWELL \$1142 PWELL NAND3_X1
X$744 \$3 NWELL PWELL FILLCELL_X8
X$745 \$3 NWELL PWELL FILLCELL_X4
X$746 \$1222 \$3 NWELL \$1101 PWELL CLKBUF_X1
X$747 \$1253 \$1254 \$3 NWELL \$772 PWELL NAND2_X1
X$748 \$3 NWELL PWELL FILLCELL_X4
X$749 \$3 NWELL PWELL NWELL TAPCELL_X1
X$750 \$3 NWELL PWELL FILLCELL_X1
X$751 \$3 NWELL PWELL FILLCELL_X2
X$752 \$123 \$999 \$3 NWELL \$366 PWELL OR2_X2
X$753 \$690 b[2] \$3 NWELL \$914 PWELL OR2_X1
X$754 \$3 NWELL PWELL FILLCELL_X1
X$755 \$3 NWELL PWELL FILLCELL_X2
X$756 \$227 \$1050 \$3 NWELL \$1157 PWELL NOR2_X1
X$757 \$914 \$3 NWELL \$1088 PWELL CLKBUF_X1
X$758 \$3 NWELL PWELL FILLCELL_X1
X$759 \$3 NWELL PWELL FILLCELL_X4
X$760 \$3 NWELL PWELL FILLCELL_X2
X$761 \$366 \$3 NWELL \$335 PWELL INV_X1
X$762 \$3 NWELL PWELL FILLCELL_X2
X$763 \$1178 \$913 \$1108 \$3 \$1089 NWELL PWELL AOI21_X1
X$764 \$3 NWELL PWELL FILLCELL_X4
X$765 \$3 NWELL PWELL FILLCELL_X4
X$766 \$1108 \$913 \$909 NWELL \$551 \$3 PWELL OAI21_X1
X$767 \$3 NWELL PWELL FILLCELL_X2
X$768 \$3 NWELL PWELL FILLCELL_X1
X$769 \$913 \$1177 \$1182 NWELL \$3 \$919 PWELL OAI21_X2
X$770 \$1242 \$3 NWELL \$1109 PWELL CLKBUF_X1
X$771 \$917 \$1001 \$1182 \$3 NWELL \$1153 PWELL NAND3_X1
X$772 \$3 NWELL PWELL FILLCELL_X1
X$773 \$3 NWELL PWELL FILLCELL_X4
X$774 \$3 NWELL PWELL FILLCELL_X2
X$775 \$3 NWELL PWELL FILLCELL_X2
X$776 \$3 NWELL PWELL FILLCELL_X1
X$777 \$1157 \$3 NWELL \$1111 PWELL CLKBUF_X1
X$778 \$3 NWELL PWELL FILLCELL_X2
X$779 NWELL VIA_via1_2_940_340_1_3_300_300
X$780 NWELL VIA_via2_3_940_340_1_3_320_320
X$781 NWELL VIA_via3_4_940_340_1_3_320_320
X$782 NWELL VIA_via1_2_940_340_1_3_300_300
X$783 NWELL VIA_via2_3_940_340_1_3_320_320
X$784 NWELL VIA_via3_4_940_340_1_3_320_320
X$785 \$3 NWELL PWELL FILLCELL_X8
X$786 \$3 NWELL PWELL NWELL TAPCELL_X1
X$787 a[2] \$3 NWELL \$690 PWELL CLKBUF_X1
X$788 a[2] \$200 NWELL \$3 \$534 PWELL AND2_X1
X$789 \$279 \$606 \$645 NWELL \$474 \$3 PWELL OAI21_X1
X$790 \$534 a[1] \$90 \$3 \$354 NWELL PWELL AOI21_X2
X$791 \$3 NWELL PWELL FILLCELL_X2
X$792 \$3 NWELL PWELL NWELL TAPCELL_X1
X$793 a[0] \$3 NWELL \$1162 PWELL CLKBUF_X1
X$794 \$3 NWELL PWELL FILLCELL_X4
X$795 \$3 NWELL PWELL FILLCELL_X2
X$796 \$3 NWELL PWELL FILLCELL_X1
X$797 b[2] \$3 NWELL \$818 PWELL CLKBUF_X1
X$798 \$3 NWELL PWELL FILLCELL_X32
X$799 NWELL VIA_via1_2_940_340_1_3_300_300
X$800 NWELL VIA_via2_3_940_340_1_3_320_320
X$801 NWELL VIA_via3_4_940_340_1_3_320_320
X$802 \$3 NWELL PWELL FILLCELL_X2
X$803 \$801 \$173 \$354 NWELL \$3 \$230 PWELL OAI21_X2
X$804 \$3 NWELL PWELL FILLCELL_X32
X$805 \$174 \$574 \$612 NWELL \$794 \$3 PWELL OAI21_X1
X$806 \$3 NWELL PWELL FILLCELL_X4
X$807 \$3 NWELL PWELL NWELL TAPCELL_X1
X$808 \$3 NWELL PWELL FILLCELL_X16
X$809 \$3 NWELL PWELL FILLCELL_X2
X$810 \$3 NWELL PWELL FILLCELL_X8
X$811 \$3 NWELL PWELL FILLCELL_X1
X$812 \$769 \$289 \$614 \$770 \$3 \$819 NWELL PWELL AOI211_X1
X$813 \$769 \$825 \$772 \$606 \$3 NWELL \$599 PWELL OR4_X1
X$814 \$769 \$770 \$289 \$3 NWELL \$960 PWELL OR3_X1
X$815 NWELL VIA_via1_2_940_340_1_3_300_300
X$816 NWELL VIA_via2_3_940_340_1_3_320_320
X$817 NWELL VIA_via3_4_940_340_1_3_320_320
X$818 \$772 \$825 \$3 NWELL \$231 PWELL NOR2_X1
X$819 \$827 \$3 NWELL \$360 PWELL CLKBUF_X1
X$820 \$3 NWELL PWELL FILLCELL_X16
X$821 \$3 NWELL PWELL FILLCELL_X8
X$822 \$723 \$3 NWELL \$711 PWELL CLKBUF_X1
X$823 \$3 NWELL PWELL FILLCELL_X1
X$824 \$619 \$3 NWELL \$620 PWELL CLKBUF_X1
X$825 \$709 \$3 NWELL \$708 PWELL CLKBUF_X1
X$826 \$620 \$3 NWELL \$723 PWELL INV_X1
X$827 \$3 NWELL PWELL FILLCELL_X1
X$828 \$593 \$3 NWELL \$809 PWELL CLKBUF_X1
X$829 \$3 NWELL PWELL FILLCELL_X8
X$830 \$3 NWELL PWELL FILLCELL_X4
X$831 \$3 NWELL PWELL FILLCELL_X2
X$832 \$3 NWELL PWELL FILLCELL_X2
X$833 \$833 \$104 \$552 \$3 NWELL \$917 PWELL NOR3_X1
X$834 \$3 NWELL PWELL FILLCELL_X2
X$835 \$3 NWELL PWELL FILLCELL_X1
X$836 \$549 \$551 NWELL \$3 \$808 PWELL XNOR2_X1
X$837 \$3 NWELL PWELL FILLCELL_X2
X$838 \$777 \$63 \$62 \$3 NWELL \$838 PWELL NOR3_X1
X$839 NWELL VIA_via1_2_940_340_1_3_300_300
X$840 NWELL VIA_via2_3_940_340_1_3_320_320
X$841 NWELL VIA_via3_4_940_340_1_3_320_320
X$842 \$879 \$838 \$809 \$3 NWELL \$980 PWELL OR3_X1
X$843 \$3 NWELL PWELL FILLCELL_X2
X$844 \$737 \$3 NWELL PWELL LOGIC0_X1
X$845 \$808 \$294 \$3 NWELL \$879 PWELL NOR2_X1
X$846 \$3 NWELL PWELL FILLCELL_X8
X$847 \$747 \$3 NWELL PWELL LOGIC0_X1
X$848 \$3 NWELL PWELL FILLCELL_X1
X$849 \$3 NWELL PWELL FILLCELL_X4
X$850 \$3 NWELL PWELL FILLCELL_X2
X$851 \$3 NWELL PWELL FILLCELL_X2
X$852 \$3 NWELL PWELL FILLCELL_X8
X$853 \$438 \$3 NWELL \$779 PWELL CLKBUF_X1
X$854 \$3 NWELL PWELL FILLCELL_X4
X$855 \$3 NWELL PWELL FILLCELL_X2
X$856 \$3 NWELL PWELL FILLCELL_X2
X$857 \$554 \$3 NWELL \$778 PWELL INV_X1
X$858 \$778 \$197 \$3 NWELL \$1003 PWELL NAND2_X1
X$859 \$3 NWELL PWELL FILLCELL_X4
X$860 \$3 NWELL PWELL FILLCELL_X2
X$861 \$779 \$427 \$780 \$839 \$3 NWELL \$866 PWELL NOR4_X1
X$862 \$779 \$3 NWELL \$862 PWELL INV_X1
X$863 \$3 NWELL PWELL FILLCELL_X1
X$864 \$3 NWELL PWELL NWELL TAPCELL_X1
X$865 \$3 NWELL PWELL FILLCELL_X4
X$866 \$555 \$3 NWELL \$753 PWELL CLKBUF_X1
X$867 \$3 NWELL PWELL FILLCELL_X1
X$868 \$3 NWELL PWELL FILLCELL_X4
X$869 \$3 NWELL PWELL FILLCELL_X2
X$870 \$3 NWELL PWELL FILLCELL_X2
X$871 \$862 \$3 NWELL \$860 PWELL CLKBUF_X1
X$872 \$840 \$3 NWELL PWELL LOGIC0_X1
X$873 \$3 NWELL PWELL FILLCELL_X1
X$874 \$957 \$557 \$780 \$3 NWELL \$843 PWELL MUX2_X1
X$875 \$744 \$3 NWELL \$735 PWELL CLKBUF_X1
X$876 \$3 NWELL PWELL FILLCELL_X1
X$877 \$747 \$3 NWELL \$758 PWELL INV_X1
X$878 \$3 NWELL PWELL FILLCELL_X2
X$879 NWELL VIA_via1_2_940_340_1_3_300_300
X$880 NWELL VIA_via2_3_940_340_1_3_320_320
X$881 NWELL VIA_via3_4_940_340_1_3_320_320
X$882 \$3 NWELL PWELL FILLCELL_X2
X$883 \$3 NWELL PWELL FILLCELL_X32
X$884 \$3 NWELL PWELL NWELL TAPCELL_X1
X$885 \$3 NWELL PWELL FILLCELL_X32
X$886 \$3 NWELL PWELL FILLCELL_X8
X$887 \$3 NWELL PWELL FILLCELL_X4
X$888 \$3 NWELL PWELL FILLCELL_X1
X$889 \$3 NWELL PWELL NWELL TAPCELL_X1
X$890 \$3 NWELL PWELL FILLCELL_X32
X$891 \$3 NWELL PWELL FILLCELL_X32
X$892 \$3 NWELL PWELL FILLCELL_X8
X$893 \$3 NWELL PWELL FILLCELL_X4
X$894 \$3 NWELL PWELL FILLCELL_X1
X$895 \$3 NWELL PWELL NWELL TAPCELL_X1
X$896 \$3 NWELL PWELL FILLCELL_X32
X$897 \$3 NWELL PWELL FILLCELL_X32
X$898 \$3 NWELL PWELL FILLCELL_X8
X$899 \$3 NWELL PWELL FILLCELL_X4
X$900 \$3 NWELL PWELL FILLCELL_X1
X$901 \$3 NWELL PWELL NWELL TAPCELL_X1
X$902 \$3 NWELL PWELL FILLCELL_X16
X$903 \$3 NWELL PWELL FILLCELL_X8
X$904 \$3 NWELL PWELL FILLCELL_X2
X$905 \$3 NWELL PWELL NWELL TAPCELL_X1
X$906 \$3 NWELL PWELL FILLCELL_X32
X$907 NWELL VIA_via1_2_940_340_1_3_300_300
X$908 NWELL VIA_via2_3_940_340_1_3_320_320
X$909 NWELL VIA_via3_4_940_340_1_3_320_320
X$910 \$3 NWELL PWELL FILLCELL_X32
X$911 \$3 NWELL PWELL FILLCELL_X32
X$912 NWELL VIA_via1_2_940_340_1_3_300_300
X$913 NWELL VIA_via2_3_940_340_1_3_320_320
X$914 NWELL VIA_via3_4_940_340_1_3_320_320
X$915 \$3 NWELL PWELL FILLCELL_X32
X$916 NWELL VIA_via1_2_940_340_1_3_300_300
X$917 NWELL VIA_via2_3_940_340_1_3_320_320
X$918 NWELL VIA_via3_4_940_340_1_3_320_320
X$919 \$3 NWELL PWELL FILLCELL_X16
X$920 \$3 NWELL PWELL FILLCELL_X8
X$921 \$3 NWELL PWELL FILLCELL_X4
X$922 \$3 NWELL PWELL NWELL TAPCELL_X1
X$923 \$3 NWELL PWELL FILLCELL_X32
X$924 NWELL VIA_via1_2_940_340_1_3_300_300
X$925 NWELL VIA_via2_3_940_340_1_3_320_320
X$926 NWELL VIA_via3_4_940_340_1_3_320_320
X$927 \$3 NWELL PWELL FILLCELL_X32
X$928 \$3 NWELL PWELL FILLCELL_X32
X$929 NWELL VIA_via1_2_940_340_1_3_300_300
X$930 NWELL VIA_via2_3_940_340_1_3_320_320
X$931 NWELL VIA_via3_4_940_340_1_3_320_320
X$932 \$3 NWELL PWELL FILLCELL_X4
X$933 \$3 NWELL PWELL FILLCELL_X2
X$934 \$3 NWELL PWELL FILLCELL_X1
X$935 \$3 NWELL PWELL NWELL TAPCELL_X1
X$936 \$3 NWELL PWELL NWELL TAPCELL_X1
X$937 \$3 NWELL PWELL NWELL TAPCELL_X1
X$938 \$3 NWELL PWELL NWELL TAPCELL_X1
X$939 \$3 NWELL PWELL FILLCELL_X32
X$940 \$3 NWELL PWELL FILLCELL_X32
X$941 NWELL VIA_via1_2_940_340_1_3_300_300
X$942 NWELL VIA_via2_3_940_340_1_3_320_320
X$943 NWELL VIA_via3_4_940_340_1_3_320_320
X$944 \$3 NWELL PWELL FILLCELL_X32
X$945 \$3 NWELL PWELL FILLCELL_X32
X$946 \$3 NWELL PWELL FILLCELL_X8
X$947 \$3 NWELL PWELL FILLCELL_X32
X$948 NWELL VIA_via1_2_940_340_1_3_300_300
X$949 NWELL VIA_via2_3_940_340_1_3_320_320
X$950 NWELL VIA_via3_4_940_340_1_3_320_320
X$951 \$3 NWELL PWELL FILLCELL_X4
X$952 \$3 NWELL PWELL FILLCELL_X1
X$953 \$3 NWELL PWELL NWELL TAPCELL_X1
X$954 \$3 NWELL PWELL FILLCELL_X32
X$955 \$3 NWELL PWELL FILLCELL_X32
X$956 \$3 NWELL PWELL FILLCELL_X32
X$957 NWELL VIA_via1_2_940_340_1_3_300_300
X$958 NWELL VIA_via2_3_940_340_1_3_320_320
X$959 NWELL VIA_via3_4_940_340_1_3_320_320
X$960 \$3 NWELL PWELL FILLCELL_X16
X$961 \$3 NWELL PWELL FILLCELL_X32
X$962 \$3 NWELL PWELL FILLCELL_X8
X$963 \$3 NWELL PWELL FILLCELL_X4
X$964 \$3 NWELL PWELL NWELL TAPCELL_X1
X$965 \$3 NWELL PWELL FILLCELL_X32
X$966 NWELL VIA_via1_2_940_340_1_3_300_300
X$967 NWELL VIA_via2_3_940_340_1_3_320_320
X$968 NWELL VIA_via3_4_940_340_1_3_320_320
X$969 \$3 NWELL PWELL FILLCELL_X32
X$970 \$3 NWELL PWELL FILLCELL_X32
X$971 \$3 NWELL PWELL FILLCELL_X16
X$972 \$3 NWELL PWELL FILLCELL_X32
X$973 \$3 NWELL PWELL FILLCELL_X8
X$974 NWELL VIA_via1_2_940_340_1_3_300_300
X$975 NWELL VIA_via2_3_940_340_1_3_320_320
X$976 NWELL VIA_via3_4_940_340_1_3_320_320
X$977 \$3 NWELL PWELL FILLCELL_X4
X$978 \$3 NWELL PWELL NWELL TAPCELL_X1
X$979 \$3 NWELL PWELL FILLCELL_X16
X$980 \$3 NWELL PWELL FILLCELL_X8
X$981 \$3 NWELL PWELL FILLCELL_X4
X$982 \$3 NWELL PWELL FILLCELL_X2
X$983 \$3 NWELL PWELL FILLCELL_X1
X$984 \$3 NWELL PWELL FILLCELL_X1
X$985 \$3 NWELL PWELL NWELL TAPCELL_X1
X$986 \$3 NWELL PWELL NWELL TAPCELL_X1
X$987 \$3 NWELL PWELL NWELL TAPCELL_X1
X$988 \$3 NWELL PWELL NWELL TAPCELL_X1
X$989 \$3 NWELL PWELL FILLCELL_X32
X$990 \$3 NWELL PWELL FILLCELL_X32
X$991 NWELL VIA_via1_2_940_340_1_3_300_300
X$992 NWELL VIA_via2_3_940_340_1_3_320_320
X$993 NWELL VIA_via3_4_940_340_1_3_320_320
X$994 \$3 NWELL PWELL FILLCELL_X32
X$995 \$3 NWELL PWELL FILLCELL_X32
X$996 \$3 NWELL PWELL FILLCELL_X8
X$997 \$3 NWELL PWELL FILLCELL_X32
X$998 NWELL VIA_via1_2_940_340_1_3_300_300
X$999 NWELL VIA_via2_3_940_340_1_3_320_320
X$1000 NWELL VIA_via3_4_940_340_1_3_320_320
X$1001 \$3 NWELL PWELL FILLCELL_X4
X$1002 \$3 NWELL PWELL FILLCELL_X1
X$1003 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1004 \$3 NWELL PWELL FILLCELL_X32
X$1005 \$3 NWELL PWELL FILLCELL_X32
X$1006 \$3 NWELL PWELL FILLCELL_X32
X$1007 NWELL VIA_via1_2_940_340_1_3_300_300
X$1008 NWELL VIA_via2_3_940_340_1_3_320_320
X$1009 NWELL VIA_via3_4_940_340_1_3_320_320
X$1010 \$3 NWELL PWELL FILLCELL_X16
X$1011 \$3 NWELL PWELL FILLCELL_X32
X$1012 \$3 NWELL PWELL FILLCELL_X8
X$1013 \$3 NWELL PWELL FILLCELL_X4
X$1014 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1015 \$3 NWELL PWELL FILLCELL_X32
X$1016 NWELL VIA_via1_2_940_340_1_3_300_300
X$1017 NWELL VIA_via2_3_940_340_1_3_320_320
X$1018 NWELL VIA_via3_4_940_340_1_3_320_320
X$1019 \$3 NWELL PWELL FILLCELL_X32
X$1020 \$3 NWELL PWELL FILLCELL_X32
X$1021 \$3 NWELL PWELL FILLCELL_X16
X$1022 \$3 NWELL PWELL FILLCELL_X32
X$1023 \$3 NWELL PWELL FILLCELL_X8
X$1024 NWELL VIA_via1_2_940_340_1_3_300_300
X$1025 NWELL VIA_via2_3_940_340_1_3_320_320
X$1026 NWELL VIA_via3_4_940_340_1_3_320_320
X$1027 \$3 NWELL PWELL FILLCELL_X4
X$1028 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1029 \$3 NWELL PWELL FILLCELL_X16
X$1030 \$3 NWELL PWELL FILLCELL_X8
X$1031 \$3 NWELL PWELL FILLCELL_X4
X$1032 \$3 NWELL PWELL FILLCELL_X2
X$1033 \$3 NWELL PWELL FILLCELL_X1
X$1034 \$3 NWELL PWELL FILLCELL_X1
X$1035 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1036 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1037 \$3 NWELL PWELL FILLCELL_X32
X$1038 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1039 \$3 NWELL PWELL FILLCELL_X32
X$1040 \$3 NWELL PWELL FILLCELL_X8
X$1041 \$3 NWELL PWELL FILLCELL_X4
X$1042 \$3 NWELL PWELL FILLCELL_X1
X$1043 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1044 \$3 NWELL PWELL FILLCELL_X32
X$1045 \$3 NWELL PWELL FILLCELL_X32
X$1046 \$3 NWELL PWELL FILLCELL_X32
X$1047 \$3 NWELL PWELL FILLCELL_X32
X$1048 \$3 NWELL PWELL FILLCELL_X16
X$1049 \$3 NWELL PWELL FILLCELL_X8
X$1050 \$3 NWELL PWELL FILLCELL_X4
X$1051 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1052 \$3 NWELL PWELL FILLCELL_X16
X$1053 \$3 NWELL PWELL FILLCELL_X8
X$1054 \$3 NWELL PWELL FILLCELL_X1
X$1055 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1056 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1057 \$3 NWELL PWELL FILLCELL_X32
X$1058 NWELL VIA_via1_2_940_340_1_3_300_300
X$1059 NWELL VIA_via2_3_940_340_1_3_320_320
X$1060 NWELL VIA_via3_4_940_340_1_3_320_320
X$1061 \$3 NWELL PWELL FILLCELL_X32
X$1062 \$3 NWELL PWELL FILLCELL_X32
X$1063 NWELL VIA_via1_2_940_340_1_3_300_300
X$1064 NWELL VIA_via2_3_940_340_1_3_320_320
X$1065 NWELL VIA_via3_4_940_340_1_3_320_320
X$1066 \$3 NWELL PWELL FILLCELL_X32
X$1067 NWELL VIA_via1_2_940_340_1_3_300_300
X$1068 NWELL VIA_via2_3_940_340_1_3_320_320
X$1069 NWELL VIA_via3_4_940_340_1_3_320_320
X$1070 \$3 NWELL PWELL FILLCELL_X16
X$1071 \$3 NWELL PWELL FILLCELL_X8
X$1072 \$3 NWELL PWELL FILLCELL_X4
X$1073 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1074 \$3 NWELL PWELL FILLCELL_X32
X$1075 NWELL VIA_via1_2_940_340_1_3_300_300
X$1076 NWELL VIA_via2_3_940_340_1_3_320_320
X$1077 NWELL VIA_via3_4_940_340_1_3_320_320
X$1078 \$3 NWELL PWELL FILLCELL_X32
X$1079 \$3 NWELL PWELL FILLCELL_X32
X$1080 NWELL VIA_via1_2_940_340_1_3_300_300
X$1081 NWELL VIA_via2_3_940_340_1_3_320_320
X$1082 NWELL VIA_via3_4_940_340_1_3_320_320
X$1083 \$3 NWELL PWELL FILLCELL_X4
X$1084 \$3 NWELL PWELL FILLCELL_X2
X$1085 \$3 NWELL PWELL FILLCELL_X1
X$1086 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1087 \$3 NWELL PWELL FILLCELL_X32
X$1088 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1089 \$3 NWELL PWELL FILLCELL_X2
X$1090 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1091 \$3 NWELL PWELL FILLCELL_X16
X$1092 \$3 NWELL PWELL FILLCELL_X8
X$1093 \$3 NWELL PWELL FILLCELL_X1
X$1094 a[5] \$3 NWELL \$27 PWELL CLKBUF_X1
X$1095 \$215 \$173 \$3 NWELL \$195 PWELL NAND2_X1
X$1096 \$3 NWELL PWELL FILLCELL_X8
X$1097 \$91 \$90 a[6] \$3 \$149 NWELL PWELL AOI21_X2
X$1098 \$91 \$90 \$18 \$3 \$306 NWELL PWELL AOI21_X2
X$1099 a[6] \$90 \$27 \$3 NWELL \$127 PWELL MUX2_X1
X$1100 \$55 \$67 \$3 NWELL \$91 PWELL NOR2_X1
X$1101 \$3 NWELL PWELL FILLCELL_X2
X$1102 \$173 \$90 a[6] \$3 \$172 NWELL PWELL AOI21_X1
X$1103 \$3 NWELL PWELL FILLCELL_X1
X$1104 \$173 \$127 \$255 \$195 NWELL \$207 \$3 PWELL OAI211_X1
X$1105 \$3 NWELL PWELL FILLCELL_X2
X$1106 \$3 NWELL PWELL FILLCELL_X1
X$1107 \$197 \$174 \$200 \$3 NWELL \$128 PWELL NAND3_X1
X$1108 \$3 NWELL PWELL FILLCELL_X16
X$1109 \$3 NWELL PWELL FILLCELL_X4
X$1110 \$75 \$67 \$3 NWELL \$129 PWELL NOR2_X1
X$1111 \$17 \$55 \$3 NWELL \$56 PWELL NOR2_X1
X$1112 \$101 \$75 \$3 NWELL \$179 PWELL NOR2_X1
X$1113 a[6] \$101 \$3 NWELL \$134 PWELL OR2_X1
X$1114 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1115 \$123 \$227 \$17 \$55 \$225 NWELL \$3 PWELL AOI211_X2
X$1116 \$101 \$131 \$3 NWELL \$103 PWELL NAND2_X2
X$1117 \$134 \$103 NWELL \$3 \$206 PWELL AND2_X1
X$1118 \$3 NWELL PWELL FILLCELL_X16
X$1119 \$3 NWELL PWELL FILLCELL_X2
X$1120 \$3 NWELL PWELL FILLCELL_X4
X$1121 \$3 NWELL PWELL FILLCELL_X2
X$1122 \$3 NWELL PWELL FILLCELL_X1
X$1123 \$123 \$227 \$176 \$3 NWELL PWELL NOR2_X4
X$1124 \$265 \$207 \$203 \$3 NWELL \$132 PWELL NAND3_X1
X$1125 \$3 NWELL PWELL FILLCELL_X2
X$1126 \$3 NWELL PWELL FILLCELL_X1
X$1127 \$206 \$3 NWELL \$104 PWELL BUF_X2
X$1128 \$3 NWELL PWELL FILLCELL_X8
X$1129 \$3 NWELL PWELL FILLCELL_X4
X$1130 \$217 b[4] \$176 NWELL \$138 \$3 PWELL OAI21_X1
X$1131 \$20 \$47 \$3 NWELL \$61 PWELL NOR2_X1
X$1132 \$3 NWELL PWELL FILLCELL_X1
X$1133 \$63 \$61 \$81 \$3 NWELL \$237 PWELL OR3_X1
X$1134 \$3 NWELL PWELL FILLCELL_X1
X$1135 \$118 \$3 NWELL \$105 PWELL CLKBUF_X1
X$1136 \$3 NWELL PWELL FILLCELL_X8
X$1137 \$3 NWELL PWELL FILLCELL_X2
X$1138 \$3 NWELL PWELL FILLCELL_X1
X$1139 \$179 \$3 NWELL \$187 PWELL CLKBUF_X1
X$1140 b[4] \$18 \$3 NWELL \$180 PWELL NAND2_X1
X$1141 \$3 NWELL PWELL FILLCELL_X4
X$1142 \$56 \$183 \$26 \$3 \$186 NWELL PWELL AOI21_X1
X$1143 \$3 NWELL PWELL FILLCELL_X4
X$1144 \$103 \$134 \$3 NWELL \$185 PWELL NAND2_X1
X$1145 \$185 \$186 \$3 NWELL \$240 PWELL OR2_X1
X$1146 \$104 \$105 \$44 \$3 \$141 NWELL PWELL AOI21_X2
X$1147 \$3 NWELL PWELL FILLCELL_X1
X$1148 \$105 \$44 \$104 \$3 NWELL \$143 PWELL NAND3_X1
X$1149 \$143 \$3 NWELL \$142 PWELL CLKBUF_X1
X$1150 \$63 \$141 \$3 NWELL \$144 PWELL NOR2_X1
X$1151 \$3 NWELL PWELL FILLCELL_X32
X$1152 \$3 NWELL PWELL FILLCELL_X32
X$1153 \$3 NWELL PWELL FILLCELL_X8
X$1154 \$3 NWELL PWELL FILLCELL_X4
X$1155 \$3 NWELL PWELL FILLCELL_X2
X$1156 \$141 \$179 \$238 NWELL \$295 \$3 PWELL OAI21_X1
X$1157 \$144 \$142 \$132 \$242 \$240 \$245 NWELL \$3 PWELL AOI221_X2
X$1158 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1159 \$141 \$187 \$3 NWELL \$374 PWELL NOR2_X1
X$1160 \$3 NWELL PWELL FILLCELL_X32
X$1161 \$3 NWELL PWELL FILLCELL_X32
X$1162 \$3 NWELL PWELL FILLCELL_X32
X$1163 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1164 \$3 NWELL PWELL FILLCELL_X1
X$1165 \$3 NWELL PWELL FILLCELL_X16
X$1166 \$3 NWELL PWELL FILLCELL_X8
X$1167 \$3 NWELL PWELL FILLCELL_X1
X$1168 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1169 \$3 NWELL PWELL FILLCELL_X4
X$1170 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1171 NWELL VIA_via1_2_940_340_1_3_300_300
X$1172 NWELL VIA_via2_3_940_340_1_3_320_320
X$1173 NWELL VIA_via3_4_940_340_1_3_320_320
X$1174 NWELL VIA_via1_2_940_340_1_3_300_300
X$1175 NWELL VIA_via2_3_940_340_1_3_320_320
X$1176 NWELL VIA_via3_4_940_340_1_3_320_320
X$1177 NWELL VIA_via1_2_940_340_1_3_300_300
X$1178 NWELL VIA_via2_3_940_340_1_3_320_320
X$1179 NWELL VIA_via3_4_940_340_1_3_320_320
X$1180 NWELL VIA_via1_2_940_340_1_3_300_300
X$1181 NWELL VIA_via2_3_940_340_1_3_320_320
X$1182 NWELL VIA_via3_4_940_340_1_3_320_320
X$1183 NWELL VIA_via1_2_940_340_1_3_300_300
X$1184 NWELL VIA_via2_3_940_340_1_3_320_320
X$1185 NWELL VIA_via3_4_940_340_1_3_320_320
X$1186 \$3 NWELL PWELL FILLCELL_X32
X$1187 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1188 \$3 NWELL PWELL FILLCELL_X32
X$1189 \$3 NWELL PWELL FILLCELL_X8
X$1190 \$3 NWELL PWELL FILLCELL_X4
X$1191 \$3 NWELL PWELL FILLCELL_X1
X$1192 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1193 \$3 NWELL PWELL FILLCELL_X32
X$1194 \$3 NWELL PWELL FILLCELL_X32
X$1195 \$3 NWELL PWELL FILLCELL_X32
X$1196 \$3 NWELL PWELL FILLCELL_X32
X$1197 \$3 NWELL PWELL FILLCELL_X16
X$1198 \$3 NWELL PWELL FILLCELL_X8
X$1199 \$3 NWELL PWELL FILLCELL_X4
X$1200 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1201 \$3 NWELL PWELL FILLCELL_X16
X$1202 \$3 NWELL PWELL FILLCELL_X8
X$1203 \$3 NWELL PWELL FILLCELL_X1
X$1204 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1205 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1206 \$3 NWELL PWELL FILLCELL_X32
X$1207 NWELL VIA_via1_2_940_340_1_3_300_300
X$1208 NWELL VIA_via2_3_940_340_1_3_320_320
X$1209 NWELL VIA_via3_4_940_340_1_3_320_320
X$1210 \$3 NWELL PWELL FILLCELL_X32
X$1211 \$3 NWELL PWELL FILLCELL_X32
X$1212 NWELL VIA_via1_2_940_340_1_3_300_300
X$1213 NWELL VIA_via2_3_940_340_1_3_320_320
X$1214 NWELL VIA_via3_4_940_340_1_3_320_320
X$1215 \$3 NWELL PWELL FILLCELL_X32
X$1216 NWELL VIA_via1_2_940_340_1_3_300_300
X$1217 NWELL VIA_via2_3_940_340_1_3_320_320
X$1218 NWELL VIA_via3_4_940_340_1_3_320_320
X$1219 \$3 NWELL PWELL FILLCELL_X16
X$1220 \$3 NWELL PWELL FILLCELL_X8
X$1221 \$3 NWELL PWELL FILLCELL_X4
X$1222 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1223 \$3 NWELL PWELL FILLCELL_X32
X$1224 NWELL VIA_via1_2_940_340_1_3_300_300
X$1225 NWELL VIA_via2_3_940_340_1_3_320_320
X$1226 NWELL VIA_via3_4_940_340_1_3_320_320
X$1227 \$3 NWELL PWELL FILLCELL_X32
X$1228 \$3 NWELL PWELL FILLCELL_X32
X$1229 NWELL VIA_via1_2_940_340_1_3_300_300
X$1230 NWELL VIA_via2_3_940_340_1_3_320_320
X$1231 NWELL VIA_via3_4_940_340_1_3_320_320
X$1232 \$3 NWELL PWELL FILLCELL_X4
X$1233 \$3 NWELL PWELL FILLCELL_X2
X$1234 \$3 NWELL PWELL FILLCELL_X1
X$1235 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1236 \$3 NWELL PWELL FILLCELL_X32
X$1237 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1238 \$3 NWELL PWELL FILLCELL_X16
X$1239 \$3 NWELL PWELL FILLCELL_X8
X$1240 \$3 NWELL PWELL FILLCELL_X4
X$1241 \$3 NWELL PWELL FILLCELL_X1
X$1242 \$1314 \$1338 \$3 \$123 NWELL PWELL OR2_X4
X$1243 \$3 NWELL PWELL FILLCELL_X4
X$1244 \$3 NWELL PWELL FILLCELL_X2
X$1245 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1246 \$3 NWELL PWELL FILLCELL_X32
X$1247 NWELL VIA_via1_2_940_340_1_3_300_300
X$1248 NWELL VIA_via2_3_940_340_1_3_320_320
X$1249 NWELL VIA_via3_4_940_340_1_3_320_320
X$1250 \$3 NWELL PWELL FILLCELL_X16
X$1251 \$3 NWELL PWELL FILLCELL_X8
X$1252 \$3 NWELL PWELL FILLCELL_X4
X$1253 \$3 NWELL PWELL FILLCELL_X2
X$1254 \$1314 \$1315 \$3 \$998 NWELL PWELL NAND2_X4
X$1255 NWELL VIA_via1_2_940_340_1_3_300_300
X$1256 NWELL VIA_via2_3_940_340_1_3_320_320
X$1257 NWELL VIA_via3_4_940_340_1_3_320_320
X$1258 opcode[3] \$3 NWELL \$1315 PWELL INV_X1
X$1259 \$3 NWELL PWELL FILLCELL_X32
X$1260 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1261 \$3 NWELL PWELL FILLCELL_X1
X$1262 \$998 \$3 NWELL \$1050 PWELL CLKBUF_X1
X$1263 \$3 NWELL PWELL FILLCELL_X32
X$1264 \$3 NWELL PWELL FILLCELL_X32
X$1265 \$3 NWELL PWELL FILLCELL_X16
X$1266 \$1319 \$3 NWELL \$1320 PWELL CLKBUF_X1
X$1267 \$3 NWELL PWELL FILLCELL_X4
X$1268 \$3 NWELL PWELL FILLCELL_X32
X$1269 NWELL VIA_via1_2_940_340_1_3_300_300
X$1270 NWELL VIA_via2_3_940_340_1_3_320_320
X$1271 NWELL VIA_via3_4_940_340_1_3_320_320
X$1272 \$3 NWELL PWELL FILLCELL_X16
X$1273 \$3 NWELL PWELL FILLCELL_X2
X$1274 \$3 NWELL PWELL FILLCELL_X1
X$1275 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1276 \$3 NWELL PWELL FILLCELL_X32
X$1277 NWELL VIA_via1_2_940_340_1_3_300_300
X$1278 NWELL VIA_via2_3_940_340_1_3_320_320
X$1279 NWELL VIA_via3_4_940_340_1_3_320_320
X$1280 \$3 NWELL PWELL FILLCELL_X16
X$1281 \$3 NWELL PWELL FILLCELL_X32
X$1282 \$3 NWELL PWELL FILLCELL_X8
X$1283 \$3 NWELL PWELL FILLCELL_X4
X$1284 \$3 NWELL PWELL FILLCELL_X2
X$1285 \$3 NWELL PWELL FILLCELL_X32
X$1286 \$3 NWELL PWELL FILLCELL_X32
X$1287 NWELL VIA_via1_2_940_340_1_3_300_300
X$1288 NWELL VIA_via2_3_940_340_1_3_320_320
X$1289 NWELL VIA_via3_4_940_340_1_3_320_320
X$1290 \$3 NWELL PWELL FILLCELL_X16
X$1291 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1292 \$3 NWELL PWELL FILLCELL_X8
X$1293 \$3 NWELL PWELL FILLCELL_X1
X$1294 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1295 \$3 NWELL PWELL FILLCELL_X4
X$1296 \$3 NWELL PWELL FILLCELL_X2
X$1297 \$3 NWELL PWELL FILLCELL_X1
X$1298 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1299 \$3 NWELL PWELL FILLCELL_X32
X$1300 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1301 \$3 NWELL PWELL FILLCELL_X32
X$1302 \$3 NWELL PWELL FILLCELL_X8
X$1303 \$3 NWELL PWELL FILLCELL_X4
X$1304 \$3 NWELL PWELL FILLCELL_X1
X$1305 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1306 \$3 NWELL PWELL FILLCELL_X32
X$1307 \$3 NWELL PWELL FILLCELL_X32
X$1308 \$3 NWELL PWELL FILLCELL_X32
X$1309 \$3 NWELL PWELL FILLCELL_X32
X$1310 \$3 NWELL PWELL FILLCELL_X16
X$1311 \$3 NWELL PWELL FILLCELL_X8
X$1312 \$3 NWELL PWELL FILLCELL_X4
X$1313 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1314 \$3 NWELL PWELL FILLCELL_X16
X$1315 \$3 NWELL PWELL FILLCELL_X8
X$1316 \$3 NWELL PWELL FILLCELL_X1
X$1317 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1318 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1319 \$3 NWELL PWELL FILLCELL_X32
X$1320 NWELL VIA_via1_2_940_340_1_3_300_300
X$1321 \$3 NWELL PWELL FILLCELL_X32
X$1322 \$3 NWELL PWELL FILLCELL_X32
X$1323 NWELL VIA_via1_2_940_340_1_3_300_300
X$1324 \$3 NWELL PWELL FILLCELL_X32
X$1325 NWELL VIA_via1_2_940_340_1_3_300_300
X$1326 \$3 NWELL PWELL FILLCELL_X16
X$1327 \$3 NWELL PWELL FILLCELL_X8
X$1328 \$3 NWELL PWELL FILLCELL_X4
X$1329 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1330 \$3 NWELL PWELL FILLCELL_X32
X$1331 NWELL VIA_via1_2_940_340_1_3_300_300
X$1332 \$3 NWELL PWELL FILLCELL_X32
X$1333 \$3 NWELL PWELL FILLCELL_X32
X$1334 NWELL VIA_via1_2_940_340_1_3_300_300
X$1335 \$3 NWELL PWELL FILLCELL_X4
X$1336 \$3 NWELL PWELL FILLCELL_X2
X$1337 \$3 NWELL PWELL FILLCELL_X1
X$1338 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1339 NWELL VIA_via2_3_940_340_1_3_320_320
X$1340 NWELL VIA_via3_4_940_340_1_3_320_320
X$1341 NWELL VIA_via2_3_940_340_1_3_320_320
X$1342 NWELL VIA_via3_4_940_340_1_3_320_320
X$1343 NWELL VIA_via2_3_940_340_1_3_320_320
X$1344 NWELL VIA_via3_4_940_340_1_3_320_320
X$1345 NWELL VIA_via2_3_940_340_1_3_320_320
X$1346 NWELL VIA_via3_4_940_340_1_3_320_320
X$1347 NWELL VIA_via2_3_940_340_1_3_320_320
X$1348 NWELL VIA_via3_4_940_340_1_3_320_320
X$1349 \$3 NWELL PWELL FILLCELL_X32
X$1350 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1351 \$3 NWELL PWELL FILLCELL_X32
X$1352 \$3 NWELL PWELL FILLCELL_X8
X$1353 \$3 NWELL PWELL FILLCELL_X4
X$1354 \$3 NWELL PWELL FILLCELL_X1
X$1355 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1356 \$3 NWELL PWELL FILLCELL_X32
X$1357 \$3 NWELL PWELL FILLCELL_X32
X$1358 \$3 NWELL PWELL FILLCELL_X32
X$1359 \$3 NWELL PWELL FILLCELL_X32
X$1360 \$3 NWELL PWELL FILLCELL_X16
X$1361 \$3 NWELL PWELL FILLCELL_X8
X$1362 \$3 NWELL PWELL FILLCELL_X4
X$1363 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1364 \$3 NWELL PWELL FILLCELL_X16
X$1365 \$3 NWELL PWELL FILLCELL_X8
X$1366 \$3 NWELL PWELL FILLCELL_X1
X$1367 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1368 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1369 \$3 NWELL PWELL FILLCELL_X32
X$1370 NWELL VIA_via1_2_940_340_1_3_300_300
X$1371 NWELL VIA_via2_3_940_340_1_3_320_320
X$1372 NWELL VIA_via3_4_940_340_1_3_320_320
X$1373 \$3 NWELL PWELL FILLCELL_X32
X$1374 \$3 NWELL PWELL FILLCELL_X16
X$1375 NWELL VIA_via1_2_940_340_1_3_300_300
X$1376 NWELL VIA_via2_3_940_340_1_3_320_320
X$1377 NWELL VIA_via3_4_940_340_1_3_320_320
X$1378 \$3 NWELL PWELL FILLCELL_X8
X$1379 \$3 NWELL PWELL FILLCELL_X4
X$1380 b[5] \$3 NWELL \$17 PWELL INV_X1
X$1381 \$3 NWELL PWELL FILLCELL_X8
X$1382 \$3 NWELL PWELL FILLCELL_X4
X$1383 \$3 NWELL PWELL FILLCELL_X1
X$1384 b[4] \$18 NWELL \$20 \$3 PWELL XOR2_X2
X$1385 \$3 NWELL PWELL FILLCELL_X1
X$1386 \$34 \$18 \$3 NWELL \$23 PWELL NAND2_X1
X$1387 NWELL VIA_via1_2_940_340_1_3_300_300
X$1388 NWELL VIA_via2_3_940_340_1_3_320_320
X$1389 NWELL VIA_via3_4_940_340_1_3_320_320
X$1390 \$3 NWELL PWELL FILLCELL_X32
X$1391 \$3 NWELL PWELL FILLCELL_X4
X$1392 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1393 \$3 NWELL PWELL FILLCELL_X32
X$1394 NWELL VIA_via1_2_940_340_1_3_300_300
X$1395 NWELL VIA_via2_3_940_340_1_3_320_320
X$1396 NWELL VIA_via3_4_940_340_1_3_320_320
X$1397 \$3 NWELL PWELL FILLCELL_X32
X$1398 \$3 NWELL PWELL FILLCELL_X32
X$1399 NWELL VIA_via1_2_940_340_1_3_300_300
X$1400 NWELL VIA_via2_3_940_340_1_3_320_320
X$1401 NWELL VIA_via3_4_940_340_1_3_320_320
X$1402 \$3 NWELL PWELL FILLCELL_X4
X$1403 \$3 NWELL PWELL FILLCELL_X2
X$1404 \$3 NWELL PWELL FILLCELL_X1
X$1405 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1406 \$3 NWELL PWELL FILLCELL_X32
X$1407 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1408 \$3 NWELL PWELL FILLCELL_X32
X$1409 \$3 NWELL PWELL FILLCELL_X8
X$1410 \$3 NWELL PWELL FILLCELL_X4
X$1411 \$3 NWELL PWELL FILLCELL_X1
X$1412 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1413 \$3 NWELL PWELL FILLCELL_X32
X$1414 \$3 NWELL PWELL FILLCELL_X32
X$1415 \$3 NWELL PWELL FILLCELL_X32
X$1416 \$3 NWELL PWELL FILLCELL_X32
X$1417 \$3 NWELL PWELL FILLCELL_X16
X$1418 \$3 NWELL PWELL FILLCELL_X8
X$1419 \$3 NWELL PWELL FILLCELL_X4
X$1420 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1421 \$3 NWELL PWELL FILLCELL_X16
X$1422 \$3 NWELL PWELL FILLCELL_X8
X$1423 \$3 NWELL PWELL FILLCELL_X1
X$1424 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1425 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1426 \$3 NWELL PWELL FILLCELL_X32
X$1427 NWELL VIA_via1_2_940_340_1_3_300_300
X$1428 NWELL VIA_via2_3_940_340_1_3_320_320
X$1429 NWELL VIA_via3_4_940_340_1_3_320_320
X$1430 \$3 NWELL PWELL FILLCELL_X32
X$1431 \$3 NWELL PWELL FILLCELL_X8
X$1432 NWELL VIA_via1_2_940_340_1_3_300_300
X$1433 NWELL VIA_via2_3_940_340_1_3_320_320
X$1434 NWELL VIA_via3_4_940_340_1_3_320_320
X$1435 \$3 NWELL PWELL FILLCELL_X4
X$1436 \$3 NWELL PWELL FILLCELL_X1
X$1437 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1438 \$3 NWELL PWELL FILLCELL_X8
X$1439 \$3 NWELL PWELL FILLCELL_X4
X$1440 \$3 NWELL PWELL FILLCELL_X2
X$1441 \$3 NWELL PWELL FILLCELL_X1
X$1442 opcode[0] \$3 NWELL \$1305 PWELL CLKBUF_X1
X$1443 opcode[3] \$3 NWELL \$1338 PWELL CLKBUF_X1
X$1444 opcode[2] \$3 NWELL \$1314 PWELL CLKBUF_X1
X$1445 \$3 NWELL PWELL FILLCELL_X8
X$1446 \$3 NWELL PWELL FILLCELL_X1
X$1447 opcode[0] \$3 NWELL \$1254 PWELL CLKBUF_X1
X$1448 \$3 NWELL PWELL FILLCELL_X32
X$1449 NWELL VIA_via1_2_940_340_1_3_300_300
X$1450 NWELL VIA_via2_3_940_340_1_3_320_320
X$1451 NWELL VIA_via3_4_940_340_1_3_320_320
X$1452 \$3 NWELL PWELL FILLCELL_X8
X$1453 \$3 NWELL PWELL FILLCELL_X1
X$1454 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1455 \$3 NWELL PWELL FILLCELL_X32
X$1456 NWELL VIA_via1_2_940_340_1_3_300_300
X$1457 NWELL VIA_via2_3_940_340_1_3_320_320
X$1458 NWELL VIA_via3_4_940_340_1_3_320_320
X$1459 \$3 NWELL PWELL FILLCELL_X32
X$1460 \$3 NWELL PWELL FILLCELL_X8
X$1461 NWELL VIA_via1_2_940_340_1_3_300_300
X$1462 NWELL VIA_via2_3_940_340_1_3_320_320
X$1463 NWELL VIA_via3_4_940_340_1_3_320_320
X$1464 \$3 NWELL PWELL FILLCELL_X4
X$1465 \$3 NWELL PWELL FILLCELL_X1
X$1466 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1467 \$3 NWELL PWELL FILLCELL_X16
X$1468 \$3 NWELL PWELL FILLCELL_X8
X$1469 \$3 NWELL PWELL FILLCELL_X2
X$1470 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1471 \$3 NWELL PWELL FILLCELL_X32
X$1472 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1473 \$3 NWELL PWELL FILLCELL_X32
X$1474 \$3 NWELL PWELL FILLCELL_X8
X$1475 \$3 NWELL PWELL FILLCELL_X4
X$1476 \$3 NWELL PWELL FILLCELL_X1
X$1477 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1478 \$3 NWELL PWELL FILLCELL_X4
X$1479 \$3 NWELL PWELL FILLCELL_X2
X$1480 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1481 \$3 NWELL PWELL FILLCELL_X32
X$1482 \$3 NWELL PWELL FILLCELL_X8
X$1483 \$18 \$67 a[5] \$3 NWELL \$126 PWELL MUX2_X1
X$1484 \$3 NWELL PWELL FILLCELL_X8
X$1485 \$3 NWELL PWELL FILLCELL_X4
X$1486 \$27 \$3 NWELL \$55 PWELL INV_X1
X$1487 \$3 NWELL PWELL FILLCELL_X4
X$1488 \$3 NWELL PWELL FILLCELL_X2
X$1489 a[6] \$3 NWELL \$75 PWELL INV_X1
X$1490 \$3 NWELL PWELL FILLCELL_X16
X$1491 b[5] \$27 NWELL \$26 \$3 PWELL XOR2_X2
X$1492 \$27 b[5] \$3 NWELL \$40 PWELL XNOR2_X2
X$1493 \$3 NWELL PWELL FILLCELL_X4
X$1494 \$3 NWELL PWELL FILLCELL_X2
X$1495 \$3 NWELL PWELL FILLCELL_X8
X$1496 \$3 NWELL PWELL FILLCELL_X4
X$1497 \$3 NWELL PWELL FILLCELL_X2
X$1498 \$3 NWELL PWELL FILLCELL_X1
X$1499 \$31 \$27 \$17 \$3 \$118 NWELL PWELL AOI21_X2
X$1500 \$3 NWELL PWELL FILLCELL_X1
X$1501 \$30 \$40 \$3 NWELL \$162 PWELL NAND2_X1
X$1502 \$3 NWELL PWELL FILLCELL_X4
X$1503 \$18 b[4] \$3 NWELL \$30 PWELL XNOR2_X2
X$1504 \$3 NWELL PWELL FILLCELL_X1
X$1505 b[4] \$3 NWELL \$34 PWELL INV_X1
X$1506 \$23 \$26 \$3 NWELL \$43 PWELL NAND2_X1
X$1507 \$23 \$26 \$3 NWELL \$31 PWELL NOR2_X1
X$1508 \$3 NWELL PWELL FILLCELL_X32
X$1509 \$3 NWELL PWELL FILLCELL_X32
X$1510 \$3 NWELL PWELL FILLCELL_X32
X$1511 \$3 NWELL PWELL FILLCELL_X4
X$1512 \$3 NWELL PWELL FILLCELL_X2
X$1513 \$30 \$62 \$42 \$3 NWELL \$81 PWELL NOR3_X1
X$1514 \$40 \$30 \$62 \$42 \$44 \$3 NWELL PWELL OAI211_X2
X$1515 \$61 \$43 \$44 \$45 NWELL \$72 \$3 PWELL OAI211_X1
X$1516 \$63 \$31 \$3 NWELL \$45 PWELL NOR2_X1
X$1517 \$62 \$42 \$3 NWELL \$47 PWELL NOR2_X1
X$1518 \$3 NWELL PWELL FILLCELL_X16
X$1519 \$3 NWELL PWELL FILLCELL_X4
X$1520 \$3 NWELL PWELL FILLCELL_X1
X$1521 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1522 \$3 NWELL PWELL FILLCELL_X32
X$1523 \$3 NWELL PWELL FILLCELL_X32
X$1524 \$3 NWELL PWELL FILLCELL_X32
X$1525 \$3 NWELL PWELL FILLCELL_X16
X$1526 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1527 \$3 NWELL PWELL FILLCELL_X8
X$1528 \$3 NWELL PWELL FILLCELL_X1
X$1529 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1530 \$3 NWELL PWELL FILLCELL_X4
X$1531 \$3 NWELL PWELL FILLCELL_X2
X$1532 \$3 NWELL PWELL FILLCELL_X1
X$1533 \$3 NWELL PWELL NWELL TAPCELL_X1
X$1534 NWELL VIA_via1_2_940_340_1_3_300_300
X$1535 NWELL VIA_via2_3_940_340_1_3_320_320
X$1536 NWELL VIA_via3_4_940_340_1_3_320_320
X$1537 NWELL VIA_via1_2_940_340_1_3_300_300
X$1538 NWELL VIA_via2_3_940_340_1_3_320_320
X$1539 NWELL VIA_via3_4_940_340_1_3_320_320
X$1540 NWELL VIA_via1_2_940_340_1_3_300_300
X$1541 NWELL VIA_via2_3_940_340_1_3_320_320
X$1542 NWELL VIA_via3_4_940_340_1_3_320_320
X$1543 NWELL VIA_via1_2_940_340_1_3_300_300
X$1544 NWELL VIA_via2_3_940_340_1_3_320_320
X$1545 NWELL VIA_via3_4_940_340_1_3_320_320
X$1546 NWELL VIA_via1_2_940_340_1_3_300_300
X$1547 NWELL VIA_via2_3_940_340_1_3_320_320
X$1548 NWELL VIA_via3_4_940_340_1_3_320_320
X$1549 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1550 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1551 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1552 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1553 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1554 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1555 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1556 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1557 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1558 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1559 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1560 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1561 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1562 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1563 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1564 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1565 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1566 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1567 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1568 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1569 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1570 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1571 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1572 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1573 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1574 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1575 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1576 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1577 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1578 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1579 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1580 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1581 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1582 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1583 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1584 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1585 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1586 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1587 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1588 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1589 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1590 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1591 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1592 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1593 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1594 NWELL VIA_via5_6_940_1600_3_2_600_600
X$1595 NWELL VIA_via4_5_940_1600_3_2_600_600
X$1596 NWELL VIA_via6_7_940_1600_2_1_600_600
X$1597 NWELL VIA_via7_8_940_1600_1_1_1680_1680
X$1598 NWELL VIA_via8_9_940_1600_1_1_1680_1680
X$1599 \$3 VIA_via9_10_1600_1600_1_1_3360_3360
X$1600 \$3 VIA_via9_10_1600_1600_1_1_3360_3360
X$1601 \$3 VIA_via9_10_1600_1600_1_1_3360_3360
X$1602 \$3 VIA_via9_10_1600_1600_1_1_3360_3360
X$1603 \$3 VIA_via1_2_940_340_1_3_300_300
X$1604 \$3 VIA_via2_3_940_340_1_3_320_320
X$1605 \$3 VIA_via3_4_940_340_1_3_320_320
X$1606 \$3 VIA_via1_2_940_340_1_3_300_300
X$1607 \$3 VIA_via2_3_940_340_1_3_320_320
X$1608 \$3 VIA_via3_4_940_340_1_3_320_320
X$1609 \$3 VIA_via1_2_940_340_1_3_300_300
X$1610 \$3 VIA_via2_3_940_340_1_3_320_320
X$1611 \$3 VIA_via3_4_940_340_1_3_320_320
X$1612 \$3 VIA_via1_2_940_340_1_3_300_300
X$1613 \$3 VIA_via2_3_940_340_1_3_320_320
X$1614 \$3 VIA_via3_4_940_340_1_3_320_320
X$1615 \$3 VIA_via1_2_940_340_1_3_300_300
X$1616 \$3 VIA_via2_3_940_340_1_3_320_320
X$1617 \$3 VIA_via3_4_940_340_1_3_320_320
X$1618 \$3 VIA_via1_2_940_340_1_3_300_300
X$1619 \$3 VIA_via2_3_940_340_1_3_320_320
X$1620 \$3 VIA_via3_4_940_340_1_3_320_320
X$1621 \$3 VIA_via1_2_940_340_1_3_300_300
X$1622 \$3 VIA_via2_3_940_340_1_3_320_320
X$1623 \$3 VIA_via3_4_940_340_1_3_320_320
X$1624 \$3 VIA_via1_2_940_340_1_3_300_300
X$1625 \$3 VIA_via2_3_940_340_1_3_320_320
X$1626 \$3 VIA_via3_4_940_340_1_3_320_320
X$1627 \$3 VIA_via1_2_940_340_1_3_300_300
X$1628 \$3 VIA_via2_3_940_340_1_3_320_320
X$1629 \$3 VIA_via3_4_940_340_1_3_320_320
X$1630 \$3 VIA_via1_2_940_340_1_3_300_300
X$1631 \$3 VIA_via2_3_940_340_1_3_320_320
X$1632 \$3 VIA_via3_4_940_340_1_3_320_320
X$1633 \$3 VIA_via1_2_940_340_1_3_300_300
X$1634 \$3 VIA_via2_3_940_340_1_3_320_320
X$1635 \$3 VIA_via3_4_940_340_1_3_320_320
X$1636 \$3 VIA_via1_2_940_340_1_3_300_300
X$1637 \$3 VIA_via2_3_940_340_1_3_320_320
X$1638 \$3 VIA_via3_4_940_340_1_3_320_320
X$1639 \$3 VIA_via1_2_940_340_1_3_300_300
X$1640 \$3 VIA_via2_3_940_340_1_3_320_320
X$1641 \$3 VIA_via3_4_940_340_1_3_320_320
X$1642 \$3 VIA_via1_2_940_340_1_3_300_300
X$1643 \$3 VIA_via2_3_940_340_1_3_320_320
X$1644 \$3 VIA_via3_4_940_340_1_3_320_320
X$1645 \$3 VIA_via1_2_940_340_1_3_300_300
X$1646 \$3 VIA_via2_3_940_340_1_3_320_320
X$1647 \$3 VIA_via3_4_940_340_1_3_320_320
X$1648 \$3 VIA_via1_2_940_340_1_3_300_300
X$1649 \$3 VIA_via2_3_940_340_1_3_320_320
X$1650 \$3 VIA_via3_4_940_340_1_3_320_320
X$1651 \$3 VIA_via1_2_940_340_1_3_300_300
X$1652 \$3 VIA_via2_3_940_340_1_3_320_320
X$1653 \$3 VIA_via3_4_940_340_1_3_320_320
X$1654 \$3 VIA_via1_2_940_340_1_3_300_300
X$1655 \$3 VIA_via2_3_940_340_1_3_320_320
X$1656 \$3 VIA_via3_4_940_340_1_3_320_320
X$1657 \$3 VIA_via1_2_940_340_1_3_300_300
X$1658 \$3 VIA_via2_3_940_340_1_3_320_320
X$1659 \$3 VIA_via3_4_940_340_1_3_320_320
X$1660 \$3 VIA_via5_6_940_960_2_2_600_600
X$1661 \$3 VIA_via4_5_940_960_2_2_600_600
X$1662 \$3 VIA_via6_7_940_960_1_1_600_600
X$1663 \$3 VIA_via5_6_940_960_2_2_600_600
X$1664 \$3 VIA_via4_5_940_960_2_2_600_600
X$1665 \$3 VIA_via6_7_940_960_1_1_600_600
X$1666 \$3 VIA_via5_6_940_960_2_2_600_600
X$1667 \$3 VIA_via4_5_940_960_2_2_600_600
X$1668 \$3 VIA_via6_7_940_960_1_1_600_600
X$1669 \$3 VIA_via5_6_940_960_2_2_600_600
X$1670 \$3 VIA_via4_5_940_960_2_2_600_600
X$1671 \$3 VIA_via6_7_940_960_1_1_600_600
X$1672 \$3 VIA_via5_6_940_960_2_2_600_600
X$1673 \$3 VIA_via4_5_940_960_2_2_600_600
X$1674 \$3 VIA_via6_7_940_960_1_1_600_600
X$1675 \$3 VIA_via5_6_940_960_2_2_600_600
X$1676 \$3 VIA_via4_5_940_960_2_2_600_600
X$1677 \$3 VIA_via6_7_940_960_1_1_600_600
X$1678 \$3 VIA_via5_6_940_960_2_2_600_600
X$1679 \$3 VIA_via4_5_940_960_2_2_600_600
X$1680 \$3 VIA_via6_7_940_960_1_1_600_600
X$1681 \$3 VIA_via5_6_940_960_2_2_600_600
X$1682 \$3 VIA_via4_5_940_960_2_2_600_600
X$1683 \$3 VIA_via6_7_940_960_1_1_600_600
X$1684 \$3 VIA_via5_6_940_960_2_2_600_600
X$1685 \$3 VIA_via4_5_940_960_2_2_600_600
X$1686 \$3 VIA_via6_7_940_960_1_1_600_600
X$1687 \$3 VIA_via5_6_940_960_2_2_600_600
X$1688 \$3 VIA_via4_5_940_960_2_2_600_600
X$1689 \$3 VIA_via6_7_940_960_1_1_600_600
X$1690 \$3 VIA_via5_6_940_960_2_2_600_600
X$1691 \$3 VIA_via4_5_940_960_2_2_600_600
X$1692 \$3 VIA_via6_7_940_960_1_1_600_600
X$1693 \$3 VIA_via5_6_940_960_2_2_600_600
X$1694 \$3 VIA_via4_5_940_960_2_2_600_600
X$1695 \$3 VIA_via6_7_940_960_1_1_600_600
X$1696 \$3 VIA_via5_6_940_960_2_2_600_600
X$1697 \$3 VIA_via4_5_940_960_2_2_600_600
X$1698 \$3 VIA_via6_7_940_960_1_1_600_600
X$1699 \$3 VIA_via5_6_940_960_2_2_600_600
X$1700 \$3 VIA_via4_5_940_960_2_2_600_600
X$1701 \$3 VIA_via6_7_940_960_1_1_600_600
X$1702 \$3 VIA_via5_6_940_960_2_2_600_600
X$1703 \$3 VIA_via4_5_940_960_2_2_600_600
X$1704 \$3 VIA_via6_7_940_960_1_1_600_600
X$1705 \$3 VIA_via5_6_940_960_2_2_600_600
X$1706 \$3 VIA_via4_5_940_960_2_2_600_600
X$1707 \$3 VIA_via6_7_940_960_1_1_600_600
X$1708 \$3 VIA_via5_6_940_960_2_2_600_600
X$1709 \$3 VIA_via4_5_940_960_2_2_600_600
X$1710 \$3 VIA_via6_7_940_960_1_1_600_600
X$1711 \$3 VIA_via5_6_940_960_2_2_600_600
X$1712 \$3 VIA_via4_5_940_960_2_2_600_600
X$1713 \$3 VIA_via6_7_940_960_1_1_600_600
X$1714 \$3 VIA_via5_6_940_960_2_2_600_600
X$1715 \$3 VIA_via4_5_940_960_2_2_600_600
X$1716 \$3 VIA_via6_7_940_960_1_1_600_600
X$1717 \$3 VIA_via5_6_940_960_2_2_600_600
X$1718 \$3 VIA_via4_5_940_960_2_2_600_600
X$1719 \$3 VIA_via6_7_940_960_1_1_600_600
X$1720 \$3 VIA_via5_6_940_960_2_2_600_600
X$1721 \$3 VIA_via4_5_940_960_2_2_600_600
X$1722 \$3 VIA_via6_7_940_960_1_1_600_600
X$1723 \$3 VIA_via5_6_940_960_2_2_600_600
X$1724 \$3 VIA_via4_5_940_960_2_2_600_600
X$1725 \$3 VIA_via6_7_940_960_1_1_600_600
X$1726 \$3 VIA_via5_6_940_960_2_2_600_600
X$1727 \$3 VIA_via4_5_940_960_2_2_600_600
X$1728 \$3 VIA_via6_7_940_960_1_1_600_600
X$1729 \$3 VIA_via5_6_940_960_2_2_600_600
X$1730 \$3 VIA_via4_5_940_960_2_2_600_600
X$1731 \$3 VIA_via6_7_940_960_1_1_600_600
X$1732 \$3 VIA_via5_6_940_960_2_2_600_600
X$1733 \$3 VIA_via4_5_940_960_2_2_600_600
X$1734 \$3 VIA_via6_7_940_960_1_1_600_600
X$1735 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1736 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1737 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1738 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1739 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1740 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1741 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1742 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1743 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1744 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1745 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1746 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1747 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1748 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1749 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1750 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1751 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1752 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1753 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1754 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1755 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1756 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1757 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1758 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1759 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1760 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1761 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1762 \$3 VIA_via9_10_1600_2400_1_1_3360_3360
X$1763 \$3 VIA_via8_9_1600_1600_1_1_1680_1680
X$1764 \$3 VIA_via7_8_1600_960_1_1_1680_1680
X$1765 \$3 VIA_via1_2_940_340_1_3_300_300
X$1766 \$3 VIA_via2_3_940_340_1_3_320_320
X$1767 \$3 VIA_via3_4_940_340_1_3_320_320
X$1768 \$3 VIA_via1_2_940_340_1_3_300_300
X$1769 \$3 VIA_via2_3_940_340_1_3_320_320
X$1770 \$3 VIA_via3_4_940_340_1_3_320_320
X$1771 \$3 VIA_via1_2_940_340_1_3_300_300
X$1772 \$3 VIA_via2_3_940_340_1_3_320_320
X$1773 \$3 VIA_via3_4_940_340_1_3_320_320
X$1774 \$3 VIA_via1_2_940_340_1_3_300_300
X$1775 \$3 VIA_via2_3_940_340_1_3_320_320
X$1776 \$3 VIA_via3_4_940_340_1_3_320_320
X$1777 \$3 VIA_via1_2_940_340_1_3_300_300
X$1778 \$3 VIA_via2_3_940_340_1_3_320_320
X$1779 \$3 VIA_via3_4_940_340_1_3_320_320
X$1780 \$3 VIA_via1_2_940_340_1_3_300_300
X$1781 \$3 VIA_via2_3_940_340_1_3_320_320
X$1782 \$3 VIA_via3_4_940_340_1_3_320_320
X$1783 \$3 VIA_via1_2_940_340_1_3_300_300
X$1784 \$3 VIA_via2_3_940_340_1_3_320_320
X$1785 \$3 VIA_via3_4_940_340_1_3_320_320
X$1786 \$3 VIA_via1_2_940_340_1_3_300_300
X$1787 \$3 VIA_via2_3_940_340_1_3_320_320
X$1788 \$3 VIA_via3_4_940_340_1_3_320_320
X$1789 \$3 VIA_via1_2_940_340_1_3_300_300
X$1790 \$3 VIA_via2_3_940_340_1_3_320_320
X$1791 \$3 VIA_via3_4_940_340_1_3_320_320
X$1792 \$3 VIA_via1_2_940_340_1_3_300_300
X$1793 \$3 VIA_via2_3_940_340_1_3_320_320
X$1794 \$3 VIA_via3_4_940_340_1_3_320_320
X$1795 \$3 VIA_via1_2_940_340_1_3_300_300
X$1796 \$3 VIA_via2_3_940_340_1_3_320_320
X$1797 \$3 VIA_via3_4_940_340_1_3_320_320
X$1798 \$3 VIA_via1_2_940_340_1_3_300_300
X$1799 \$3 VIA_via2_3_940_340_1_3_320_320
X$1800 \$3 VIA_via3_4_940_340_1_3_320_320
X$1801 \$3 VIA_via1_2_940_340_1_3_300_300
X$1802 \$3 VIA_via2_3_940_340_1_3_320_320
X$1803 \$3 VIA_via3_4_940_340_1_3_320_320
X$1804 \$3 VIA_via1_2_940_340_1_3_300_300
X$1805 \$3 VIA_via2_3_940_340_1_3_320_320
X$1806 \$3 VIA_via3_4_940_340_1_3_320_320
X$1807 \$3 VIA_via1_2_940_340_1_3_300_300
X$1808 \$3 VIA_via2_3_940_340_1_3_320_320
X$1809 \$3 VIA_via3_4_940_340_1_3_320_320
X$1810 \$3 VIA_via1_2_940_340_1_3_300_300
X$1811 \$3 VIA_via2_3_940_340_1_3_320_320
X$1812 \$3 VIA_via3_4_940_340_1_3_320_320
X$1813 \$3 VIA_via1_2_940_340_1_3_300_300
X$1814 \$3 VIA_via2_3_940_340_1_3_320_320
X$1815 \$3 VIA_via3_4_940_340_1_3_320_320
X$1816 \$3 VIA_via1_2_940_340_1_3_300_300
X$1817 \$3 VIA_via2_3_940_340_1_3_320_320
X$1818 \$3 VIA_via3_4_940_340_1_3_320_320
X$1819 \$3 VIA_via1_2_940_340_1_3_300_300
X$1820 \$3 VIA_via2_3_940_340_1_3_320_320
X$1821 \$3 VIA_via3_4_940_340_1_3_320_320
X$1822 \$3 VIA_via1_2_940_340_1_3_300_300
X$1823 \$3 VIA_via2_3_940_340_1_3_320_320
X$1824 \$3 VIA_via3_4_940_340_1_3_320_320
X$1825 \$3 VIA_via1_2_940_340_1_3_300_300
X$1826 \$3 VIA_via2_3_940_340_1_3_320_320
X$1827 \$3 VIA_via3_4_940_340_1_3_320_320
X$1828 \$3 VIA_via1_2_940_340_1_3_300_300
X$1829 \$3 VIA_via2_3_940_340_1_3_320_320
X$1830 \$3 VIA_via3_4_940_340_1_3_320_320
X$1831 \$3 VIA_via1_2_940_340_1_3_300_300
X$1832 \$3 VIA_via2_3_940_340_1_3_320_320
X$1833 \$3 VIA_via3_4_940_340_1_3_320_320
X$1834 \$3 VIA_via1_2_940_340_1_3_300_300
X$1835 \$3 VIA_via2_3_940_340_1_3_320_320
X$1836 \$3 VIA_via3_4_940_340_1_3_320_320
X$1837 \$3 VIA_via1_2_940_340_1_3_300_300
X$1838 \$3 VIA_via2_3_940_340_1_3_320_320
X$1839 \$3 VIA_via3_4_940_340_1_3_320_320
X$1840 \$3 VIA_via1_2_940_340_1_3_300_300
X$1841 \$3 VIA_via2_3_940_340_1_3_320_320
X$1842 \$3 VIA_via3_4_940_340_1_3_320_320
X$1843 \$3 VIA_via1_2_940_340_1_3_300_300
X$1844 \$3 VIA_via2_3_940_340_1_3_320_320
X$1845 \$3 VIA_via3_4_940_340_1_3_320_320
X$1846 \$3 VIA_via1_2_940_340_1_3_300_300
X$1847 \$3 VIA_via2_3_940_340_1_3_320_320
X$1848 \$3 VIA_via3_4_940_340_1_3_320_320
X$1849 \$3 VIA_via1_2_940_340_1_3_300_300
X$1850 \$3 VIA_via2_3_940_340_1_3_320_320
X$1851 \$3 VIA_via3_4_940_340_1_3_320_320
X$1852 \$3 VIA_via1_2_940_340_1_3_300_300
X$1853 \$3 VIA_via2_3_940_340_1_3_320_320
X$1854 \$3 VIA_via3_4_940_340_1_3_320_320
X$1855 \$3 VIA_via1_2_940_340_1_3_300_300
X$1856 \$3 VIA_via2_3_940_340_1_3_320_320
X$1857 \$3 VIA_via3_4_940_340_1_3_320_320
X$1858 \$3 VIA_via1_2_940_340_1_3_300_300
X$1859 \$3 VIA_via2_3_940_340_1_3_320_320
X$1860 \$3 VIA_via3_4_940_340_1_3_320_320
X$1861 \$3 VIA_via1_2_940_340_1_3_300_300
X$1862 \$3 VIA_via2_3_940_340_1_3_320_320
X$1863 \$3 VIA_via3_4_940_340_1_3_320_320
X$1864 \$3 VIA_via1_2_940_340_1_3_300_300
X$1865 \$3 VIA_via2_3_940_340_1_3_320_320
X$1866 \$3 VIA_via3_4_940_340_1_3_320_320
X$1867 \$3 VIA_via1_2_940_340_1_3_300_300
X$1868 \$3 VIA_via2_3_940_340_1_3_320_320
X$1869 \$3 VIA_via3_4_940_340_1_3_320_320
X$1870 \$3 VIA_via1_2_940_340_1_3_300_300
X$1871 \$3 VIA_via2_3_940_340_1_3_320_320
X$1872 \$3 VIA_via3_4_940_340_1_3_320_320
X$1873 \$3 VIA_via1_2_940_340_1_3_300_300
X$1874 \$3 VIA_via2_3_940_340_1_3_320_320
X$1875 \$3 VIA_via3_4_940_340_1_3_320_320
X$1876 \$3 VIA_via1_2_940_340_1_3_300_300
X$1877 \$3 VIA_via2_3_940_340_1_3_320_320
X$1878 \$3 VIA_via3_4_940_340_1_3_320_320
X$1879 \$3 VIA_via1_2_940_340_1_3_300_300
X$1880 \$3 VIA_via2_3_940_340_1_3_320_320
X$1881 \$3 VIA_via3_4_940_340_1_3_320_320
X$1882 \$3 VIA_via1_2_940_340_1_3_300_300
X$1883 \$3 VIA_via2_3_940_340_1_3_320_320
X$1884 \$3 VIA_via3_4_940_340_1_3_320_320
X$1885 \$3 VIA_via1_2_940_340_1_3_300_300
X$1886 \$3 VIA_via2_3_940_340_1_3_320_320
X$1887 \$3 VIA_via3_4_940_340_1_3_320_320
X$1888 \$3 VIA_via1_2_940_340_1_3_300_300
X$1889 \$3 VIA_via2_3_940_340_1_3_320_320
X$1890 \$3 VIA_via3_4_940_340_1_3_320_320
X$1891 \$3 VIA_via1_2_940_340_1_3_300_300
X$1892 \$3 VIA_via2_3_940_340_1_3_320_320
X$1893 \$3 VIA_via3_4_940_340_1_3_320_320
X$1894 \$3 VIA_via1_2_940_340_1_3_300_300
X$1895 \$3 VIA_via2_3_940_340_1_3_320_320
X$1896 \$3 VIA_via3_4_940_340_1_3_320_320
X$1897 \$3 VIA_via1_2_940_340_1_3_300_300
X$1898 \$3 VIA_via2_3_940_340_1_3_320_320
X$1899 \$3 VIA_via3_4_940_340_1_3_320_320
X$1900 \$3 VIA_via1_2_940_340_1_3_300_300
X$1901 \$3 VIA_via2_3_940_340_1_3_320_320
X$1902 \$3 VIA_via3_4_940_340_1_3_320_320
X$1903 \$3 VIA_via1_2_940_340_1_3_300_300
X$1904 \$3 VIA_via2_3_940_340_1_3_320_320
X$1905 \$3 VIA_via3_4_940_340_1_3_320_320
X$1906 \$3 VIA_via1_2_940_340_1_3_300_300
X$1907 \$3 VIA_via2_3_940_340_1_3_320_320
X$1908 \$3 VIA_via3_4_940_340_1_3_320_320
X$1909 \$3 VIA_via1_2_940_340_1_3_300_300
X$1910 \$3 VIA_via2_3_940_340_1_3_320_320
X$1911 \$3 VIA_via3_4_940_340_1_3_320_320
X$1912 \$3 VIA_via1_2_940_340_1_3_300_300
X$1913 \$3 VIA_via2_3_940_340_1_3_320_320
X$1914 \$3 VIA_via3_4_940_340_1_3_320_320
X$1915 \$3 VIA_via1_2_940_340_1_3_300_300
X$1916 \$3 VIA_via2_3_940_340_1_3_320_320
X$1917 \$3 VIA_via3_4_940_340_1_3_320_320
X$1918 \$3 VIA_via1_2_940_340_1_3_300_300
X$1919 \$3 VIA_via2_3_940_340_1_3_320_320
X$1920 \$3 VIA_via3_4_940_340_1_3_320_320
X$1921 \$3 VIA_via1_2_940_340_1_3_300_300
X$1922 \$3 VIA_via2_3_940_340_1_3_320_320
X$1923 \$3 VIA_via3_4_940_340_1_3_320_320
X$1924 \$3 VIA_via1_2_940_340_1_3_300_300
X$1925 \$3 VIA_via2_3_940_340_1_3_320_320
X$1926 \$3 VIA_via3_4_940_340_1_3_320_320
X$1927 \$3 VIA_via1_2_940_340_1_3_300_300
X$1928 \$3 VIA_via2_3_940_340_1_3_320_320
X$1929 \$3 VIA_via3_4_940_340_1_3_320_320
X$1930 \$3 VIA_via1_2_940_340_1_3_300_300
X$1931 \$3 VIA_via2_3_940_340_1_3_320_320
X$1932 \$3 VIA_via3_4_940_340_1_3_320_320
X$1933 \$3 VIA_via1_2_940_340_1_3_300_300
X$1934 \$3 VIA_via2_3_940_340_1_3_320_320
X$1935 \$3 VIA_via3_4_940_340_1_3_320_320
X$1936 \$3 VIA_via1_2_940_340_1_3_300_300
X$1937 \$3 VIA_via2_3_940_340_1_3_320_320
X$1938 \$3 VIA_via3_4_940_340_1_3_320_320
X$1939 \$3 VIA_via1_2_940_340_1_3_300_300
X$1940 \$3 VIA_via2_3_940_340_1_3_320_320
X$1941 \$3 VIA_via3_4_940_340_1_3_320_320
X$1942 \$3 VIA_via1_2_940_340_1_3_300_300
X$1943 \$3 VIA_via2_3_940_340_1_3_320_320
X$1944 \$3 VIA_via3_4_940_340_1_3_320_320
X$1945 \$3 VIA_via1_2_940_340_1_3_300_300
X$1946 \$3 VIA_via2_3_940_340_1_3_320_320
X$1947 \$3 VIA_via3_4_940_340_1_3_320_320
X$1948 \$3 VIA_via1_2_940_340_1_3_300_300
X$1949 \$3 VIA_via2_3_940_340_1_3_320_320
X$1950 \$3 VIA_via3_4_940_340_1_3_320_320
X$1951 \$3 VIA_via1_2_940_340_1_3_300_300
X$1952 \$3 VIA_via2_3_940_340_1_3_320_320
X$1953 \$3 VIA_via3_4_940_340_1_3_320_320
X$1954 \$3 VIA_via1_2_940_340_1_3_300_300
X$1955 \$3 VIA_via2_3_940_340_1_3_320_320
X$1956 \$3 VIA_via3_4_940_340_1_3_320_320
X$1957 \$3 VIA_via1_2_940_340_1_3_300_300
X$1958 \$3 VIA_via2_3_940_340_1_3_320_320
X$1959 \$3 VIA_via3_4_940_340_1_3_320_320
X$1960 \$3 VIA_via1_2_940_340_1_3_300_300
X$1961 \$3 VIA_via2_3_940_340_1_3_320_320
X$1962 \$3 VIA_via3_4_940_340_1_3_320_320
X$1963 \$3 VIA_via1_2_940_340_1_3_300_300
X$1964 \$3 VIA_via2_3_940_340_1_3_320_320
X$1965 \$3 VIA_via3_4_940_340_1_3_320_320
X$1966 \$3 VIA_via1_2_940_340_1_3_300_300
X$1967 \$3 VIA_via2_3_940_340_1_3_320_320
X$1968 \$3 VIA_via3_4_940_340_1_3_320_320
X$1969 \$3 VIA_via1_2_940_340_1_3_300_300
X$1970 \$3 VIA_via2_3_940_340_1_3_320_320
X$1971 \$3 VIA_via3_4_940_340_1_3_320_320
X$1972 \$3 VIA_via1_2_940_340_1_3_300_300
X$1973 \$3 VIA_via2_3_940_340_1_3_320_320
X$1974 \$3 VIA_via3_4_940_340_1_3_320_320
X$1975 \$3 VIA_via1_2_940_340_1_3_300_300
X$1976 \$3 VIA_via2_3_940_340_1_3_320_320
X$1977 \$3 VIA_via3_4_940_340_1_3_320_320
X$1978 \$3 VIA_via5_6_940_1600_3_2_600_600
X$1979 \$3 VIA_via4_5_940_1600_3_2_600_600
X$1980 \$3 VIA_via6_7_940_1600_2_1_600_600
X$1981 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$1982 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$1983 \$3 VIA_via5_6_940_1600_3_2_600_600
X$1984 \$3 VIA_via4_5_940_1600_3_2_600_600
X$1985 \$3 VIA_via6_7_940_1600_2_1_600_600
X$1986 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$1987 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$1988 \$3 VIA_via5_6_940_1600_3_2_600_600
X$1989 \$3 VIA_via4_5_940_1600_3_2_600_600
X$1990 \$3 VIA_via6_7_940_1600_2_1_600_600
X$1991 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$1992 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$1993 \$3 VIA_via5_6_940_1600_3_2_600_600
X$1994 \$3 VIA_via4_5_940_1600_3_2_600_600
X$1995 \$3 VIA_via6_7_940_1600_2_1_600_600
X$1996 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$1997 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$1998 \$3 VIA_via5_6_940_1600_3_2_600_600
X$1999 \$3 VIA_via4_5_940_1600_3_2_600_600
X$2000 \$3 VIA_via6_7_940_1600_2_1_600_600
X$2001 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$2002 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$2003 \$3 VIA_via5_6_940_1600_3_2_600_600
X$2004 \$3 VIA_via4_5_940_1600_3_2_600_600
X$2005 \$3 VIA_via6_7_940_1600_2_1_600_600
X$2006 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$2007 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$2008 \$3 VIA_via5_6_940_1600_3_2_600_600
X$2009 \$3 VIA_via4_5_940_1600_3_2_600_600
X$2010 \$3 VIA_via6_7_940_1600_2_1_600_600
X$2011 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$2012 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$2013 \$3 VIA_via5_6_940_1600_3_2_600_600
X$2014 \$3 VIA_via4_5_940_1600_3_2_600_600
X$2015 \$3 VIA_via6_7_940_1600_2_1_600_600
X$2016 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$2017 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$2018 \$3 VIA_via5_6_940_1600_3_2_600_600
X$2019 \$3 VIA_via4_5_940_1600_3_2_600_600
X$2020 \$3 VIA_via6_7_940_1600_2_1_600_600
X$2021 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$2022 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$2023 \$3 VIA_via5_6_940_1600_3_2_600_600
X$2024 \$3 VIA_via4_5_940_1600_3_2_600_600
X$2025 \$3 VIA_via6_7_940_1600_2_1_600_600
X$2026 \$3 VIA_via7_8_940_1600_1_1_1680_1680
X$2027 \$3 VIA_via8_9_940_1600_1_1_1680_1680
X$2028 b[5] VIA_via2_5
X$2029 b[5] VIA_via2_5
X$2030 b[5] VIA_via2_5
X$2031 b[5] VIA_via2_5
X$2032 b[5] VIA_via2_5
X$2033 b[5] VIA_via1_4
X$2034 b[5] VIA_via1_4
X$2035 b[5] VIA_via2_5
X$2036 b[5] VIA_via1_4
X$2037 b[5] VIA_via2_5
X$2038 \$17 VIA_via2_5
X$2039 \$17 VIA_via2_5
X$2040 \$17 VIA_via2_5
X$2041 \$17 VIA_via2_5
X$2042 \$17 VIA_via1_4
X$2043 \$17 VIA_via1_4
X$2044 \$17 VIA_via1_4
X$2045 \$17 VIA_via1_4
X$2046 \$18 VIA_via2_5
X$2047 \$18 VIA_via2_5
X$2048 \$18 VIA_via2_5
X$2049 \$18 VIA_via2_5
X$2050 \$18 VIA_via2_5
X$2051 \$18 VIA_via2_5
X$2052 \$18 VIA_via2_5
X$2053 \$18 VIA_via2_5
X$2054 \$18 VIA_via2_5
X$2055 \$18 VIA_via2_5
X$2056 \$18 VIA_via2_5
X$2057 \$18 VIA_via2_5
X$2058 \$18 VIA_via2_5
X$2059 \$18 VIA_via1_4
X$2060 \$18 VIA_via1_4
X$2061 \$18 VIA_via1_4
X$2062 \$18 VIA_via2_5
X$2063 \$18 VIA_via1_4
X$2064 \$18 VIA_via1_4
X$2065 \$18 VIA_via2_5
X$2066 \$18 VIA_via1_4
X$2067 \$18 VIA_via1_4
X$2068 \$18 VIA_via1_4
X$2069 \$18 VIA_via1_4
X$2070 \$20 VIA_via2_5
X$2071 \$20 VIA_via2_5
X$2072 \$20 VIA_via1_4
X$2073 \$20 VIA_via1_4
X$2074 \$20 VIA_via1_4
X$2075 \$23 VIA_via2_5
X$2076 \$23 VIA_via2_5
X$2077 \$23 VIA_via1_4
X$2078 \$23 VIA_via2_5
X$2079 \$23 VIA_via1_4
X$2080 \$23 VIA_via2_5
X$2081 \$23 VIA_via1_4
X$2082 \$26 VIA_via2_5
X$2083 \$26 VIA_via3_2
X$2084 \$26 VIA_via2_5
X$2085 \$26 VIA_via3_2
X$2086 \$26 VIA_via2_5
X$2087 \$26 VIA_via1_4
X$2088 \$26 VIA_via1_4
X$2089 \$26 VIA_via1_4
X$2090 \$26 VIA_via2_5
X$2091 \$26 VIA_via1_4
X$2092 \$26 VIA_via1_4
X$2093 \$26 VIA_via2_5
X$2094 \$26 VIA_via1_4
X$2095 \$27 VIA_via2_5
X$2096 \$27 VIA_via2_5
X$2097 \$27 VIA_via2_5
X$2098 \$27 VIA_via2_5
X$2099 \$27 VIA_via2_5
X$2100 \$27 VIA_via1_4
X$2101 \$27 VIA_via1_4
X$2102 \$27 VIA_via1_4
X$2103 \$27 VIA_via2_5
X$2104 \$27 VIA_via1_4
X$2105 \$27 VIA_via2_5
X$2106 \$27 VIA_via1_4
X$2107 \$27 VIA_via2_5
X$2108 \$27 VIA_via1_4
X$2109 b[4] VIA_via3_2
X$2110 b[4] VIA_via2_5
X$2111 b[4] VIA_via2_5
X$2112 b[4] VIA_via2_5
X$2113 b[4] VIA_via1_4
X$2114 b[4] VIA_via1_4
X$2115 b[4] VIA_via2_5
X$2116 b[4] VIA_via3_2
X$2117 b[4] VIA_via1_4
X$2118 b[4] VIA_via2_5
X$2119 b[4] VIA_via1_4
X$2120 b[4] VIA_via2_5
X$2121 b[4] VIA_via3_2
X$2122 b[4] VIA_via1_4
X$2123 \$30 VIA_via2_5
X$2124 \$30 VIA_via2_5
X$2125 \$30 VIA_via2_5
X$2126 \$30 VIA_via2_5
X$2127 \$30 VIA_via2_5
X$2128 \$30 VIA_via2_5
X$2129 \$30 VIA_via2_5
X$2130 \$30 VIA_via2_5
X$2131 \$30 VIA_via1_4
X$2132 \$30 VIA_via1_4
X$2133 \$30 VIA_via1_4
X$2134 \$30 VIA_via1_4
X$2135 \$30 VIA_via1_4
X$2136 \$30 VIA_via2_5
X$2137 \$30 VIA_via1_4
X$2138 \$31 VIA_via1_4
X$2139 \$31 VIA_via1_4
X$2140 \$31 VIA_via2_5
X$2141 \$31 VIA_via1_4
X$2142 \$31 VIA_via2_5
X$2143 \$34 VIA_via2_5
X$2144 \$34 VIA_via1_4
X$2145 \$34 VIA_via2_5
X$2146 \$34 VIA_via1_4
X$2147 a[5] VIA_via2_5
X$2148 a[5] VIA_via2_5
X$2149 a[5] VIA_via2_5
X$2150 a[5] VIA_via1_4
X$2151 a[5] VIA_via1_4
X$2152 a[6] VIA_via2_5
X$2153 a[6] VIA_via2_5
X$2154 a[6] VIA_via2_5
X$2155 a[6] VIA_via2_5
X$2156 a[6] VIA_via2_5
X$2157 a[6] VIA_via2_5
X$2158 a[6] VIA_via1_4
X$2159 a[6] VIA_via1_4
X$2160 a[6] VIA_via2_5
X$2161 a[6] VIA_via1_4
X$2162 a[6] VIA_via2_5
X$2163 a[6] VIA_via1_4
X$2164 a[6] VIA_via2_5
X$2165 a[6] VIA_via1_4
X$2166 a[6] VIA_via2_5
X$2167 a[6] VIA_via1_4
X$2168 \$40 VIA_via2_5
X$2169 \$40 VIA_via1_4
X$2170 \$40 VIA_via2_5
X$2171 \$40 VIA_via2_5
X$2172 \$40 VIA_via1_4
X$2173 \$40 VIA_via1_4
X$2174 \$40 VIA_via2_5
X$2175 \$42 VIA_via2_5
X$2176 \$42 VIA_via2_5
X$2177 \$42 VIA_via2_5
X$2178 \$42 VIA_via2_5
X$2179 \$42 VIA_via2_5
X$2180 \$42 VIA_via1_4
X$2181 \$42 VIA_via2_5
X$2182 \$42 VIA_via1_4
X$2183 \$42 VIA_via1_4
X$2184 \$42 VIA_via1_4
X$2185 \$43 VIA_via1_4
X$2186 \$43 VIA_via1_4
X$2187 \$44 VIA_via2_5
X$2188 \$44 VIA_via1_4
X$2189 \$44 VIA_via2_5
X$2190 \$44 VIA_via1_4
X$2191 \$44 VIA_via2_5
X$2192 \$44 VIA_via1_4
X$2193 \$44 VIA_via2_5
X$2194 \$44 VIA_via1_4
X$2195 \$44 VIA_via2_5
X$2196 \$45 VIA_via1_4
X$2197 \$45 VIA_via1_4
X$2198 \$47 VIA_via2_5
X$2199 \$47 VIA_via1_4
X$2200 \$47 VIA_via1_4
X$2201 \$47 VIA_via2_5
X$2202 \$55 VIA_via2_5
X$2203 \$55 VIA_via1_4
X$2204 \$55 VIA_via2_5
X$2205 \$55 VIA_via1_4
X$2206 \$55 VIA_via2_5
X$2207 \$55 VIA_via1_4
X$2208 \$55 VIA_via2_5
X$2209 \$55 VIA_via1_4
X$2210 \$56 VIA_via1_7
X$2211 \$56 VIA_via1_7
X$2212 \$56 VIA_via2_5
X$2213 \$56 VIA_via2_5
X$2214 \$56 VIA_via2_5
X$2215 \$56 VIA_via1_4
X$2216 \$56 VIA_via1_4
X$2217 \$56 VIA_via1_4
X$2218 \$61 VIA_via2_5
X$2219 \$61 VIA_via2_5
X$2220 \$61 VIA_via1_4
X$2221 \$61 VIA_via2_5
X$2222 \$61 VIA_via1_4
X$2223 \$61 VIA_via1_4
X$2224 \$62 VIA_via3_2
X$2225 \$62 VIA_via3_2
X$2226 \$62 VIA_via2_5
X$2227 \$62 VIA_via2_5
X$2228 \$62 VIA_via2_5
X$2229 \$62 VIA_via2_5
X$2230 \$62 VIA_via2_5
X$2231 \$62 VIA_via2_5
X$2232 \$62 VIA_via2_5
X$2233 \$62 VIA_via2_5
X$2234 \$62 VIA_via1_4
X$2235 \$62 VIA_via1_4
X$2236 \$62 VIA_via1_4
X$2237 \$62 VIA_via1_4
X$2238 \$62 VIA_via1_4
X$2239 \$63 VIA_via2_5
X$2240 \$63 VIA_via2_5
X$2241 \$63 VIA_via2_5
X$2242 \$63 VIA_via2_5
X$2243 \$63 VIA_via2_5
X$2244 \$63 VIA_via2_5
X$2245 \$63 VIA_via2_5
X$2246 \$63 VIA_via2_5
X$2247 \$63 VIA_via2_5
X$2248 \$63 VIA_via2_5
X$2249 \$63 VIA_via2_5
X$2250 \$63 VIA_via1_4
X$2251 \$63 VIA_via1_4
X$2252 \$63 VIA_via1_4
X$2253 \$63 VIA_via1_4
X$2254 \$63 VIA_via1_4
X$2255 \$63 VIA_via1_4
X$2256 \$63 VIA_via2_5
X$2257 \$63 VIA_via1_4
X$2258 \$63 VIA_via1_4
X$2259 \$63 VIA_via1_4
X$2260 \$63 VIA_via2_5
X$2261 \$67 VIA_via2_5
X$2262 \$67 VIA_via2_5
X$2263 \$67 VIA_via2_5
X$2264 \$67 VIA_via2_5
X$2265 \$67 VIA_via2_5
X$2266 \$67 VIA_via1_4
X$2267 \$67 VIA_via1_4
X$2268 \$67 VIA_via2_5
X$2269 \$67 VIA_via1_4
X$2270 \$67 VIA_via2_5
X$2271 \$67 VIA_via1_4
X$2272 \$67 VIA_via2_5
X$2273 \$67 VIA_via1_4
X$2274 \$72 VIA_via2_5
X$2275 \$72 VIA_via2_5
X$2276 \$72 VIA_via1_4
X$2277 \$72 VIA_via1_4
X$2278 \$75 VIA_via2_5
X$2279 \$75 VIA_via1_4
X$2280 \$75 VIA_via2_5
X$2281 \$75 VIA_via1_4
X$2282 \$75 VIA_via1_4
X$2283 \$75 VIA_via2_5
X$2284 \$81 VIA_via2_5
X$2285 \$81 VIA_via2_5
X$2286 \$81 VIA_via1_4
X$2287 \$81 VIA_via1_4
X$2288 \$90 VIA_via1_7
X$2289 \$90 VIA_via1_7
X$2290 \$90 VIA_via1_7
X$2291 \$90 VIA_via1_7
X$2292 \$90 VIA_via2_5
X$2293 \$90 VIA_via2_5
X$2294 \$90 VIA_via2_5
X$2295 \$90 VIA_via2_5
X$2296 \$90 VIA_via2_5
X$2297 \$90 VIA_via2_5
X$2298 \$90 VIA_via2_5
X$2299 \$90 VIA_via2_5
X$2300 \$90 VIA_via2_5
X$2301 \$90 VIA_via1_4
X$2302 \$90 VIA_via1_4
X$2303 \$90 VIA_via2_5
X$2304 \$90 VIA_via1_4
X$2305 \$90 VIA_via1_4
X$2306 \$90 VIA_via2_5
X$2307 \$90 VIA_via1_4
X$2308 \$90 VIA_via1_4
X$2309 \$90 VIA_via1_4
X$2310 \$90 VIA_via1_4
X$2311 \$90 VIA_via2_5
X$2312 \$91 VIA_via1_4
X$2313 \$91 VIA_via2_5
X$2314 \$91 VIA_via1_4
X$2315 \$91 VIA_via2_5
X$2316 \$91 VIA_via1_4
X$2317 \$91 VIA_via2_5
X$2318 \$101 VIA_via2_5
X$2319 \$101 VIA_via2_5
X$2320 \$101 VIA_via1_4
X$2321 \$101 VIA_via2_5
X$2322 \$101 VIA_via1_4
X$2323 \$101 VIA_via1_4
X$2324 \$101 VIA_via2_5
X$2325 \$101 VIA_via1_4
X$2326 \$101 VIA_via2_5
X$2327 \$103 VIA_via2_5
X$2328 \$103 VIA_via2_5
X$2329 \$103 VIA_via2_5
X$2330 \$103 VIA_via2_5
X$2331 \$103 VIA_via2_5
X$2332 \$103 VIA_via2_5
X$2333 \$103 VIA_via2_5
X$2334 \$103 VIA_via1_4
X$2335 \$103 VIA_via2_5
X$2336 \$103 VIA_via1_4
X$2337 \$103 VIA_via1_4
X$2338 \$103 VIA_via1_4
X$2339 \$103 VIA_via1_4
X$2340 \$103 VIA_via1_4
X$2341 \$104 VIA_via3_2
X$2342 \$104 VIA_via3_2
X$2343 \$104 VIA_via2_5
X$2344 \$104 VIA_via2_5
X$2345 \$104 VIA_via2_5
X$2346 \$104 VIA_via2_5
X$2347 \$104 VIA_via1_4
X$2348 \$104 VIA_via1_4
X$2349 \$104 VIA_via1_4
X$2350 \$104 VIA_via2_5
X$2351 \$104 VIA_via1_4
X$2352 \$104 VIA_via2_5
X$2353 \$104 VIA_via1_4
X$2354 \$104 VIA_via2_5
X$2355 \$105 VIA_via1_4
X$2356 \$105 VIA_via2_5
X$2357 \$105 VIA_via1_4
X$2358 \$105 VIA_via2_5
X$2359 \$105 VIA_via1_4
X$2360 \$105 VIA_via2_5
X$2361 \$118 VIA_via2_5
X$2362 \$118 VIA_via1_4
X$2363 \$118 VIA_via1_4
X$2364 \$118 VIA_via2_5
X$2365 \$123 VIA_via2_5
X$2366 \$123 VIA_via2_5
X$2367 \$123 VIA_via2_5
X$2368 \$123 VIA_via2_5
X$2369 \$123 VIA_via2_5
X$2370 \$123 VIA_via2_5
X$2371 \$123 VIA_via2_5
X$2372 \$123 VIA_via1_4
X$2373 \$123 VIA_via1_4
X$2374 \$123 VIA_via1_4
X$2375 \$123 VIA_via1_4
X$2376 \$123 VIA_via1_4
X$2377 \$123 VIA_via1_4
X$2378 \$123 VIA_via1_4
X$2379 \$123 VIA_via2_5
X$2380 \$126 VIA_via1_7
X$2381 \$126 VIA_via1_7
X$2382 \$126 VIA_via2_5
X$2383 \$126 VIA_via2_5
X$2384 \$126 VIA_via1_4
X$2385 \$126 VIA_via2_5
X$2386 \$126 VIA_via1_4
X$2387 \$126 VIA_via2_5
X$2388 \$126 VIA_via1_4
X$2389 \$127 VIA_via1_4
X$2390 \$127 VIA_via1_4
X$2391 \$128 VIA_via2_5
X$2392 \$128 VIA_via2_5
X$2393 \$128 VIA_via1_4
X$2394 \$128 VIA_via1_4
X$2395 \$129 VIA_via1_4
X$2396 \$129 VIA_via1_4
X$2397 \$131 VIA_via2_5
X$2398 \$131 VIA_via2_5
X$2399 \$131 VIA_via1_4
X$2400 \$131 VIA_via1_4
X$2401 \$132 VIA_via2_5
X$2402 \$132 VIA_via2_5
X$2403 \$132 VIA_via1_4
X$2404 \$132 VIA_via1_4
X$2405 \$134 VIA_via2_5
X$2406 \$134 VIA_via2_5
X$2407 \$134 VIA_via2_5
X$2408 \$134 VIA_via2_5
X$2409 \$134 VIA_via1_4
X$2410 \$134 VIA_via1_4
X$2411 \$134 VIA_via1_4
X$2412 \$134 VIA_via1_4
X$2413 \$134 VIA_via2_5
X$2414 \$138 VIA_via2_5
X$2415 \$138 VIA_via2_5
X$2416 \$138 VIA_via1_4
X$2417 \$138 VIA_via1_4
X$2418 \$141 VIA_via1_7
X$2419 \$141 VIA_via2_5
X$2420 \$141 VIA_via2_5
X$2421 \$141 VIA_via2_5
X$2422 \$141 VIA_via1_4
X$2423 \$141 VIA_via1_4
X$2424 \$141 VIA_via1_4
X$2425 \$142 VIA_via1_4
X$2426 \$142 VIA_via1_4
X$2427 \$143 VIA_via1_4
X$2428 \$143 VIA_via1_4
X$2429 \$144 VIA_via1_4
X$2430 \$144 VIA_via1_4
X$2431 \$149 VIA_via1_7
X$2432 \$149 VIA_via2_5
X$2433 \$149 VIA_via2_5
X$2434 \$149 VIA_via2_5
X$2435 \$149 VIA_via2_5
X$2436 \$149 VIA_via1_4
X$2437 \$149 VIA_via1_4
X$2438 \$162 VIA_via3_2
X$2439 \$162 VIA_via2_5
X$2440 \$162 VIA_via2_5
X$2441 \$162 VIA_via3_2
X$2442 \$162 VIA_via1_4
X$2443 \$162 VIA_via1_4
X$2444 \$172 VIA_via1_4
X$2445 \$172 VIA_via1_4
X$2446 \$173 VIA_via2_5
X$2447 \$173 VIA_via2_5
X$2448 \$173 VIA_via2_5
X$2449 \$173 VIA_via2_5
X$2450 \$173 VIA_via2_5
X$2451 \$173 VIA_via2_5
X$2452 \$173 VIA_via1_4
X$2453 \$173 VIA_via1_4
X$2454 \$173 VIA_via2_5
X$2455 \$173 VIA_via1_4
X$2456 \$173 VIA_via1_4
X$2457 \$173 VIA_via1_4
X$2458 \$173 VIA_via1_4
X$2459 \$173 VIA_via1_4
X$2460 \$173 VIA_via1_4
X$2461 \$173 VIA_via2_5
X$2462 \$173 VIA_via1_4
X$2463 \$174 VIA_via2_5
X$2464 \$174 VIA_via2_5
X$2465 \$174 VIA_via2_5
X$2466 \$174 VIA_via2_5
X$2467 \$174 VIA_via2_5
X$2468 \$174 VIA_via2_5
X$2469 \$174 VIA_via2_5
X$2470 \$174 VIA_via2_5
X$2471 \$174 VIA_via1_4
X$2472 \$174 VIA_via2_5
X$2473 \$174 VIA_via1_4
X$2474 \$174 VIA_via1_4
X$2475 \$174 VIA_via1_4
X$2476 \$174 VIA_via1_4
X$2477 \$174 VIA_via1_4
X$2478 \$174 VIA_via1_4
X$2479 \$174 VIA_via1_4
X$2480 \$174 VIA_via1_4
X$2481 \$176 VIA_via3_2
X$2482 \$176 VIA_via3_2
X$2483 \$176 VIA_via3_2
X$2484 \$176 VIA_via2_5
X$2485 \$176 VIA_via3_2
X$2486 \$176 VIA_via2_5
X$2487 \$176 VIA_via2_5
X$2488 \$176 VIA_via2_5
X$2489 \$176 VIA_via2_5
X$2490 \$176 VIA_via1_4
X$2491 \$176 VIA_via1_4
X$2492 \$176 VIA_via2_5
X$2493 \$176 VIA_via3_2
X$2494 \$176 VIA_via1_4
X$2495 \$176 VIA_via2_5
X$2496 \$176 VIA_via1_4
X$2497 \$176 VIA_via2_5
X$2498 \$176 VIA_via1_4
X$2499 \$176 VIA_via1_4
X$2500 \$176 VIA_via1_4
X$2501 \$179 VIA_via2_5
X$2502 \$179 VIA_via1_4
X$2503 \$179 VIA_via2_5
X$2504 \$179 VIA_via1_4
X$2505 \$179 VIA_via2_5
X$2506 \$179 VIA_via1_4
X$2507 \$180 VIA_via1_4
X$2508 \$180 VIA_via2_5
X$2509 \$180 VIA_via1_4
X$2510 \$180 VIA_via2_5
X$2511 \$180 VIA_via1_4
X$2512 \$183 VIA_via1_4
X$2513 \$183 VIA_via2_5
X$2514 \$183 VIA_via1_4
X$2515 \$183 VIA_via1_4
X$2516 \$183 VIA_via2_5
X$2517 \$185 VIA_via2_5
X$2518 \$185 VIA_via1_4
X$2519 \$185 VIA_via1_4
X$2520 \$185 VIA_via2_5
X$2521 \$185 VIA_via1_4
X$2522 \$186 VIA_via2_5
X$2523 \$186 VIA_via2_5
X$2524 \$186 VIA_via1_4
X$2525 \$186 VIA_via2_5
X$2526 \$186 VIA_via1_4
X$2527 \$186 VIA_via1_4
X$2528 \$186 VIA_via2_5
X$2529 \$187 VIA_via2_5
X$2530 \$187 VIA_via1_4
X$2531 \$187 VIA_via2_5
X$2532 \$187 VIA_via1_4
X$2533 \$195 VIA_via1_4
X$2534 \$195 VIA_via2_5
X$2535 \$195 VIA_via1_4
X$2536 \$195 VIA_via2_5
X$2537 \$197 VIA_via2_5
X$2538 \$197 VIA_via2_5
X$2539 \$197 VIA_via2_5
X$2540 \$197 VIA_via2_5
X$2541 \$197 VIA_via2_5
X$2542 \$197 VIA_via2_5
X$2543 \$197 VIA_via2_5
X$2544 \$197 VIA_via2_5
X$2545 \$197 VIA_via2_5
X$2546 \$197 VIA_via1_4
X$2547 \$197 VIA_via1_4
X$2548 \$197 VIA_via1_4
X$2549 \$197 VIA_via1_4
X$2550 \$197 VIA_via1_4
X$2551 \$197 VIA_via2_5
X$2552 \$197 VIA_via1_4
X$2553 \$197 VIA_via1_4
X$2554 \$197 VIA_via1_4
X$2555 \$197 VIA_via1_4
X$2556 \$197 VIA_via2_5
X$2557 \$200 VIA_via3_2
X$2558 \$200 VIA_via3_2
X$2559 \$200 VIA_via3_2
X$2560 \$200 VIA_via3_2
X$2561 \$200 VIA_via2_5
X$2562 \$200 VIA_via2_5
X$2563 \$200 VIA_via2_5
X$2564 \$200 VIA_via2_5
X$2565 \$200 VIA_via2_5
X$2566 \$200 VIA_via2_5
X$2567 \$200 VIA_via1_4
X$2568 \$200 VIA_via1_4
X$2569 \$200 VIA_via2_5
X$2570 \$200 VIA_via1_4
X$2571 \$200 VIA_via2_5
X$2572 \$200 VIA_via1_4
X$2573 \$200 VIA_via1_4
X$2574 \$200 VIA_via2_5
X$2575 \$200 VIA_via1_4
X$2576 \$200 VIA_via1_4
X$2577 \$200 VIA_via2_5
X$2578 \$203 VIA_via2_5
X$2579 \$203 VIA_via1_4
X$2580 \$203 VIA_via1_4
X$2581 \$203 VIA_via2_5
X$2582 \$206 VIA_via1_4
X$2583 \$206 VIA_via1_4
X$2584 \$207 VIA_via1_4
X$2585 \$207 VIA_via2_5
X$2586 \$207 VIA_via1_4
X$2587 \$207 VIA_via2_5
X$2588 a[1] VIA_via2_5
X$2589 a[1] VIA_via2_5
X$2590 a[1] VIA_via2_5
X$2591 a[1] VIA_via2_5
X$2592 a[1] VIA_via2_5
X$2593 a[1] VIA_via2_5
X$2594 a[1] VIA_via2_5
X$2595 a[1] VIA_via2_5
X$2596 a[1] VIA_via2_5
X$2597 a[1] VIA_via2_5
X$2598 a[1] VIA_via1_4
X$2599 a[1] VIA_via1_4
X$2600 a[1] VIA_via1_4
X$2601 a[1] VIA_via1_4
X$2602 a[1] VIA_via1_4
X$2603 a[2] VIA_via2_5
X$2604 a[2] VIA_via2_5
X$2605 a[2] VIA_via2_5
X$2606 a[2] VIA_via2_5
X$2607 a[2] VIA_via2_5
X$2608 a[2] VIA_via2_5
X$2609 a[2] VIA_via2_5
X$2610 a[2] VIA_via2_5
X$2611 a[2] VIA_via1_4
X$2612 a[2] VIA_via2_5
X$2613 a[2] VIA_via1_4
X$2614 a[2] VIA_via2_5
X$2615 a[2] VIA_via1_4
X$2616 a[2] VIA_via1_4
X$2617 a[2] VIA_via1_4
X$2618 a[2] VIA_via1_4
X$2619 a[0] VIA_via2_5
X$2620 a[0] VIA_via1_4
X$2621 \$215 VIA_via2_5
X$2622 \$215 VIA_via2_5
X$2623 \$215 VIA_via2_5
X$2624 \$215 VIA_via1_4
X$2625 \$215 VIA_via1_4
X$2626 \$215 VIA_via1_4
X$2627 \$217 VIA_via2_5
X$2628 \$217 VIA_via2_5
X$2629 \$217 VIA_via1_4
X$2630 \$217 VIA_via1_4
X$2631 \$217 VIA_via2_5
X$2632 \$217 VIA_via1_4
X$2633 \$220 VIA_via2_5
X$2634 \$220 VIA_via2_5
X$2635 \$220 VIA_via1_4
X$2636 \$220 VIA_via1_4
X$2637 \$222 VIA_via2_5
X$2638 \$222 VIA_via2_5
X$2639 \$222 VIA_via2_5
X$2640 \$222 VIA_via2_5
X$2641 \$222 VIA_via2_5
X$2642 \$222 VIA_via1_4
X$2643 \$222 VIA_via1_4
X$2644 \$222 VIA_via1_4
X$2645 \$224 VIA_via3_2
X$2646 \$224 VIA_via3_2
X$2647 \$224 VIA_via3_2
X$2648 \$224 VIA_via2_5
X$2649 \$224 VIA_via2_5
X$2650 \$224 VIA_via1_4
X$2651 \$224 VIA_via2_5
X$2652 \$224 VIA_via1_4
X$2653 \$224 VIA_via2_5
X$2654 \$224 VIA_via1_4
X$2655 \$224 VIA_via2_5
X$2656 \$224 VIA_via1_4
X$2657 \$224 VIA_via1_4
X$2658 \$225 VIA_via1_4
X$2659 \$225 VIA_via1_4
X$2660 \$227 VIA_via1_7
X$2661 \$227 VIA_via3_2
X$2662 \$227 VIA_via2_5
X$2663 \$227 VIA_via3_2
X$2664 \$227 VIA_via2_5
X$2665 \$227 VIA_via2_5
X$2666 \$227 VIA_via2_5
X$2667 \$227 VIA_via2_5
X$2668 \$227 VIA_via1_4
X$2669 \$227 VIA_via1_4
X$2670 \$227 VIA_via1_4
X$2671 \$227 VIA_via2_5
X$2672 \$227 VIA_via1_4
X$2673 \$230 VIA_via2_5
X$2674 \$230 VIA_via1_4
X$2675 \$230 VIA_via1_4
X$2676 \$230 VIA_via2_5
X$2677 \$230 VIA_via1_4
X$2678 \$231 VIA_via2_5
X$2679 \$231 VIA_via2_5
X$2680 \$231 VIA_via1_4
X$2681 \$231 VIA_via1_4
X$2682 \$231 VIA_via2_5
X$2683 \$231 VIA_via1_4
X$2684 \$231 VIA_via1_4
X$2685 \$233 VIA_via3_2
X$2686 \$233 VIA_via2_5
X$2687 \$233 VIA_via2_5
X$2688 \$233 VIA_via2_5
X$2689 \$233 VIA_via2_5
X$2690 \$233 VIA_via3_2
X$2691 \$233 VIA_via2_5
X$2692 \$233 VIA_via1_4
X$2693 \$233 VIA_via1_4
X$2694 \$233 VIA_via2_5
X$2695 \$233 VIA_via1_4
X$2696 \$233 VIA_via2_5
X$2697 \$233 VIA_via1_4
X$2698 \$233 VIA_via1_4
X$2699 \$233 VIA_via1_4
X$2700 \$233 VIA_via2_5
X$2701 \$233 VIA_via1_4
X$2702 \$233 VIA_via1_4
X$2703 \$233 VIA_via2_5
X$2704 \$233 VIA_via1_4
X$2705 \$233 VIA_via2_5
X$2706 \$237 VIA_via1_4
X$2707 \$237 VIA_via1_4
X$2708 \$238 VIA_via3_2
X$2709 \$238 VIA_via3_2
X$2710 \$238 VIA_via2_5
X$2711 \$238 VIA_via1_4
X$2712 \$238 VIA_via1_4
X$2713 \$238 VIA_via1_4
X$2714 \$238 VIA_via2_5
X$2715 \$238 VIA_via1_4
X$2716 \$238 VIA_via2_5
X$2717 \$240 VIA_via2_5
X$2718 \$240 VIA_via2_5
X$2719 \$240 VIA_via2_5
X$2720 \$240 VIA_via2_5
X$2721 \$240 VIA_via1_4
X$2722 \$240 VIA_via1_4
X$2723 \$240 VIA_via1_4
X$2724 \$240 VIA_via1_4
X$2725 \$242 VIA_via1_4
X$2726 \$242 VIA_via1_4
X$2727 \$245 VIA_via3_2
X$2728 \$245 VIA_via1_4
X$2729 \$245 VIA_via2_5
X$2730 \$245 VIA_via3_2
X$2731 \$245 VIA_via1_4
X$2732 \$245 VIA_via2_5
X$2733 \$254 VIA_via2_5
X$2734 \$254 VIA_via1_4
X$2735 \$254 VIA_via1_4
X$2736 \$254 VIA_via2_5
X$2737 \$255 VIA_via3_2
X$2738 \$255 VIA_via2_5
X$2739 \$255 VIA_via2_5
X$2740 \$255 VIA_via2_5
X$2741 \$255 VIA_via2_5
X$2742 \$255 VIA_via2_5
X$2743 \$255 VIA_via2_5
X$2744 \$255 VIA_via2_5
X$2745 \$255 VIA_via1_4
X$2746 \$255 VIA_via1_4
X$2747 \$255 VIA_via1_4
X$2748 \$255 VIA_via2_5
X$2749 \$255 VIA_via3_2
X$2750 \$255 VIA_via1_4
X$2751 \$255 VIA_via1_4
X$2752 \$258 VIA_via1_7
X$2753 \$258 VIA_via2_5
X$2754 \$258 VIA_via2_5
X$2755 \$258 VIA_via1_4
X$2756 \$265 VIA_via2_5
X$2757 \$265 VIA_via2_5
X$2758 \$265 VIA_via1_4
X$2759 \$265 VIA_via1_4
X$2760 a[4] VIA_via2_5
X$2761 a[4] VIA_via1_4
X$2762 a[3] VIA_via2_5
X$2763 a[3] VIA_via2_5
X$2764 a[3] VIA_via2_5
X$2765 a[3] VIA_via1_4
X$2766 a[3] VIA_via2_5
X$2767 a[3] VIA_via1_4
X$2768 a[3] VIA_via2_5
X$2769 a[3] VIA_via1_4
X$2770 a[3] VIA_via2_5
X$2771 \$278 VIA_via2_5
X$2772 \$278 VIA_via2_5
X$2773 \$278 VIA_via1_4
X$2774 \$278 VIA_via1_4
X$2775 \$279 VIA_via2_5
X$2776 \$279 VIA_via2_5
X$2777 \$279 VIA_via2_5
X$2778 \$279 VIA_via2_5
X$2779 \$279 VIA_via2_5
X$2780 \$279 VIA_via2_5
X$2781 \$279 VIA_via2_5
X$2782 \$279 VIA_via2_5
X$2783 \$279 VIA_via2_5
X$2784 \$279 VIA_via1_4
X$2785 \$279 VIA_via1_4
X$2786 \$279 VIA_via1_4
X$2787 \$279 VIA_via2_5
X$2788 \$279 VIA_via1_4
X$2789 \$279 VIA_via1_4
X$2790 \$279 VIA_via2_5
X$2791 \$279 VIA_via1_4
X$2792 \$279 VIA_via2_5
X$2793 \$279 VIA_via1_4
X$2794 \$279 VIA_via1_4
X$2795 \$279 VIA_via2_5
X$2796 \$279 VIA_via1_4
X$2797 \$280 VIA_via1_4
X$2798 \$280 VIA_via1_4
X$2799 \$284 VIA_via2_5
X$2800 \$284 VIA_via2_5
X$2801 \$284 VIA_via2_5
X$2802 \$284 VIA_via2_5
X$2803 \$284 VIA_via2_5
X$2804 \$284 VIA_via2_5
X$2805 \$284 VIA_via2_5
X$2806 \$284 VIA_via2_5
X$2807 \$284 VIA_via1_4
X$2808 \$284 VIA_via2_5
X$2809 \$284 VIA_via1_4
X$2810 \$284 VIA_via1_4
X$2811 \$284 VIA_via1_4
X$2812 \$284 VIA_via1_4
X$2813 \$284 VIA_via1_4
X$2814 \$284 VIA_via2_5
X$2815 \$287 VIA_via2_5
X$2816 \$287 VIA_via2_5
X$2817 \$287 VIA_via2_5
X$2818 \$287 VIA_via2_5
X$2819 \$287 VIA_via2_5
X$2820 \$287 VIA_via1_4
X$2821 \$287 VIA_via1_4
X$2822 \$287 VIA_via2_5
X$2823 \$287 VIA_via1_4
X$2824 \$289 VIA_via1_7
X$2825 \$289 VIA_via2_5
X$2826 \$289 VIA_via2_5
X$2827 \$289 VIA_via2_5
X$2828 \$289 VIA_via2_5
X$2829 \$289 VIA_via2_5
X$2830 \$289 VIA_via2_5
X$2831 \$289 VIA_via1_4
X$2832 \$289 VIA_via1_4
X$2833 \$289 VIA_via1_4
X$2834 \$289 VIA_via1_4
X$2835 \$291 VIA_via2_5
X$2836 \$291 VIA_via2_5
X$2837 \$291 VIA_via1_4
X$2838 \$291 VIA_via1_4
X$2839 \$292 VIA_via1_4
X$2840 \$292 VIA_via1_4
X$2841 \$293 VIA_via1_4
X$2842 \$293 VIA_via1_4
X$2843 \$294 VIA_via2_5
X$2844 \$294 VIA_via2_5
X$2845 \$294 VIA_via2_5
X$2846 \$294 VIA_via2_5
X$2847 \$294 VIA_via2_5
X$2848 \$294 VIA_via2_5
X$2849 \$294 VIA_via2_5
X$2850 \$294 VIA_via2_5
X$2851 \$294 VIA_via2_5
X$2852 \$294 VIA_via2_5
X$2853 \$294 VIA_via1_4
X$2854 \$294 VIA_via2_5
X$2855 \$294 VIA_via1_4
X$2856 \$294 VIA_via2_5
X$2857 \$294 VIA_via1_4
X$2858 \$294 VIA_via1_4
X$2859 \$294 VIA_via1_4
X$2860 \$294 VIA_via1_4
X$2861 \$294 VIA_via1_4
X$2862 \$295 VIA_via2_5
X$2863 \$295 VIA_via2_5
X$2864 \$295 VIA_via1_4
X$2865 \$295 VIA_via1_4
X$2866 \$295 VIA_via1_4
X$2867 \$305 VIA_via2_5
X$2868 \$305 VIA_via2_5
X$2869 \$305 VIA_via1_4
X$2870 \$305 VIA_via1_4
X$2871 \$306 VIA_via1_7
X$2872 \$306 VIA_via2_5
X$2873 \$306 VIA_via1_4
X$2874 \$306 VIA_via2_5
X$2875 \$306 VIA_via1_4
X$2876 \$313 VIA_via1_7
X$2877 \$313 VIA_via2_5
X$2878 \$313 VIA_via2_5
X$2879 \$313 VIA_via2_5
X$2880 \$313 VIA_via1_4
X$2881 \$313 VIA_via1_4
X$2882 \$321 VIA_via2_5
X$2883 \$321 VIA_via2_5
X$2884 \$321 VIA_via1_4
X$2885 \$321 VIA_via1_4
X$2886 \$324 VIA_via2_5
X$2887 \$324 VIA_via2_5
X$2888 \$324 VIA_via2_5
X$2889 \$324 VIA_via2_5
X$2890 \$324 VIA_via1_4
X$2891 \$324 VIA_via1_4
X$2892 \$325 VIA_via2_5
X$2893 \$325 VIA_via2_5
X$2894 \$325 VIA_via1_4
X$2895 \$325 VIA_via1_4
X$2896 \$326 VIA_via2_5
X$2897 \$326 VIA_via2_5
X$2898 \$326 VIA_via1_4
X$2899 \$326 VIA_via1_4
X$2900 \$335 VIA_via3_2
X$2901 \$335 VIA_via3_2
X$2902 \$335 VIA_via3_2
X$2903 \$335 VIA_via2_5
X$2904 \$335 VIA_via2_5
X$2905 \$335 VIA_via2_5
X$2906 \$335 VIA_via1_4
X$2907 \$335 VIA_via1_4
X$2908 \$335 VIA_via2_5
X$2909 \$335 VIA_via1_4
X$2910 \$335 VIA_via1_4
X$2911 \$335 VIA_via2_5
X$2912 \$339 VIA_via2_5
X$2913 \$339 VIA_via2_5
X$2914 \$339 VIA_via1_4
X$2915 \$339 VIA_via1_4
X$2916 \$342 VIA_via2_5
X$2917 \$342 VIA_via1_4
X$2918 \$342 VIA_via2_5
X$2919 \$342 VIA_via1_4
X$2920 b[0] VIA_via2_5
X$2921 b[0] VIA_via1_4
X$2922 a[7] VIA_via2_5
X$2923 a[7] VIA_via2_5
X$2924 a[7] VIA_via2_5
X$2925 a[7] VIA_via1_4
X$2926 \$351 VIA_via2_5
X$2927 \$351 VIA_via2_5
X$2928 \$351 VIA_via2_5
X$2929 \$351 VIA_via1_4
X$2930 \$351 VIA_via1_4
X$2931 \$351 VIA_via1_4
X$2932 \$352 VIA_via2_5
X$2933 \$352 VIA_via1_4
X$2934 \$352 VIA_via2_5
X$2935 \$352 VIA_via1_4
X$2936 \$352 VIA_via1_4
X$2937 \$352 VIA_via2_5
X$2938 \$354 VIA_via2_5
X$2939 \$354 VIA_via1_4
X$2940 \$354 VIA_via1_4
X$2941 \$354 VIA_via1_4
X$2942 \$354 VIA_via2_5
X$2943 \$356 VIA_via1_7
X$2944 \$356 VIA_via3_2
X$2945 \$356 VIA_via3_2
X$2946 \$356 VIA_via3_2
X$2947 \$356 VIA_via2_5
X$2948 \$356 VIA_via2_5
X$2949 \$356 VIA_via2_5
X$2950 \$356 VIA_via2_5
X$2951 \$356 VIA_via2_5
X$2952 \$356 VIA_via1_4
X$2953 \$356 VIA_via2_5
X$2954 \$356 VIA_via1_4
X$2955 \$356 VIA_via1_4
X$2956 \$356 VIA_via1_4
X$2957 \$356 VIA_via1_4
X$2958 \$357 VIA_via2_5
X$2959 \$357 VIA_via2_5
X$2960 \$357 VIA_via2_5
X$2961 \$357 VIA_via2_5
X$2962 \$357 VIA_via2_5
X$2963 \$357 VIA_via2_5
X$2964 \$357 VIA_via2_5
X$2965 \$357 VIA_via2_5
X$2966 \$357 VIA_via2_5
X$2967 \$357 VIA_via2_5
X$2968 \$357 VIA_via1_4
X$2969 \$357 VIA_via1_4
X$2970 \$357 VIA_via1_4
X$2971 \$357 VIA_via1_4
X$2972 \$357 VIA_via1_4
X$2973 \$357 VIA_via1_4
X$2974 \$359 VIA_via2_5
X$2975 \$359 VIA_via1_4
X$2976 \$359 VIA_via2_5
X$2977 \$359 VIA_via1_4
X$2978 \$360 VIA_via2_5
X$2979 \$360 VIA_via2_5
X$2980 \$360 VIA_via1_4
X$2981 \$360 VIA_via1_4
X$2982 b[3] VIA_via2_5
X$2983 b[3] VIA_via2_5
X$2984 b[3] VIA_via2_5
X$2985 b[3] VIA_via2_5
X$2986 b[3] VIA_via2_5
X$2987 b[3] VIA_via2_5
X$2988 b[3] VIA_via1_4
X$2989 b[3] VIA_via1_4
X$2990 b[3] VIA_via2_5
X$2991 b[3] VIA_via1_4
X$2992 b[3] VIA_via2_5
X$2993 \$362 VIA_via2_5
X$2994 \$362 VIA_via1_4
X$2995 \$362 VIA_via1_4
X$2996 \$362 VIA_via2_5
X$2997 \$365 VIA_via1_4
X$2998 \$365 VIA_via1_4
X$2999 \$366 VIA_via3_2
X$3000 \$366 VIA_via3_2
X$3001 \$366 VIA_via3_2
X$3002 \$366 VIA_via2_5
X$3003 \$366 VIA_via2_5
X$3004 \$366 VIA_via2_5
X$3005 \$366 VIA_via2_5
X$3006 \$366 VIA_via2_5
X$3007 \$366 VIA_via2_5
X$3008 \$366 VIA_via1_4
X$3009 \$366 VIA_via1_4
X$3010 \$366 VIA_via1_4
X$3011 \$366 VIA_via1_4
X$3012 \$366 VIA_via2_5
X$3013 \$366 VIA_via1_4
X$3014 \$366 VIA_via2_5
X$3015 \$366 VIA_via1_4
X$3016 \$366 VIA_via1_4
X$3017 \$371 VIA_via2_5
X$3018 \$371 VIA_via2_5
X$3019 \$371 VIA_via1_4
X$3020 \$371 VIA_via1_4
X$3021 \$371 VIA_via1_4
X$3022 \$371 VIA_via2_5
X$3023 \$374 VIA_via2_5
X$3024 \$374 VIA_via1_4
X$3025 \$374 VIA_via2_5
X$3026 \$374 VIA_via1_4
X$3027 \$382 VIA_via2_5
X$3028 \$382 VIA_via2_5
X$3029 \$382 VIA_via2_5
X$3030 \$382 VIA_via1_4
X$3031 \$382 VIA_via2_5
X$3032 \$382 VIA_via1_4
X$3033 \$382 VIA_via1_4
X$3034 \$390 VIA_via1_4
X$3035 \$390 VIA_via1_4
X$3036 \$394 VIA_via1_4
X$3037 \$394 VIA_via2_5
X$3038 \$394 VIA_via1_4
X$3039 \$394 VIA_via2_5
X$3040 \$396 VIA_via2_5
X$3041 \$396 VIA_via1_4
X$3042 \$396 VIA_via2_5
X$3043 \$396 VIA_via1_4
X$3044 \$397 VIA_via3_2
X$3045 \$397 VIA_via3_2
X$3046 \$397 VIA_via3_2
X$3047 \$397 VIA_via2_5
X$3048 \$397 VIA_via2_5
X$3049 \$397 VIA_via2_5
X$3050 \$397 VIA_via1_4
X$3051 \$397 VIA_via2_5
X$3052 \$397 VIA_via1_4
X$3053 \$397 VIA_via1_4
X$3054 \$397 VIA_via2_5
X$3055 \$397 VIA_via1_4
X$3056 \$397 VIA_via2_5
X$3057 b[1] VIA_via2_5
X$3058 b[1] VIA_via1_4
X$3059 b[2] VIA_via2_5
X$3060 b[2] VIA_via2_5
X$3061 b[2] VIA_via2_5
X$3062 b[2] VIA_via2_5
X$3063 b[2] VIA_via2_5
X$3064 b[2] VIA_via2_5
X$3065 b[2] VIA_via2_5
X$3066 b[2] VIA_via1_4
X$3067 b[2] VIA_via1_4
X$3068 b[2] VIA_via2_5
X$3069 b[2] VIA_via1_4
X$3070 b[2] VIA_via1_4
X$3071 b[2] VIA_via2_5
X$3072 b[2] VIA_via1_4
X$3073 b[2] VIA_via2_5
X$3074 \$416 VIA_via1_7
X$3075 \$416 VIA_via1_4
X$3076 \$421 VIA_via2_5
X$3077 \$421 VIA_via1_4
X$3078 \$421 VIA_via1_4
X$3079 \$421 VIA_via2_5
X$3080 \$427 VIA_via2_5
X$3081 \$427 VIA_via1_4
X$3082 \$427 VIA_via1_4
X$3083 \$427 VIA_via1_4
X$3084 \$427 VIA_via2_5
X$3085 \$428 VIA_via2_5
X$3086 \$428 VIA_via1_4
X$3087 \$428 VIA_via1_4
X$3088 \$428 VIA_via2_5
X$3089 \$429 VIA_via2_5
X$3090 \$429 VIA_via2_5
X$3091 \$429 VIA_via1_4
X$3092 \$429 VIA_via1_4
X$3093 \$430 VIA_via2_5
X$3094 \$430 VIA_via2_5
X$3095 \$430 VIA_via1_4
X$3096 \$430 VIA_via1_4
X$3097 \$431 VIA_via2_5
X$3098 \$431 VIA_via2_5
X$3099 \$431 VIA_via1_4
X$3100 \$431 VIA_via2_5
X$3101 \$431 VIA_via1_4
X$3102 \$431 VIA_via1_4
X$3103 \$431 VIA_via1_4
X$3104 \$431 VIA_via1_4
X$3105 \$431 VIA_via1_4
X$3106 \$431 VIA_via1_4
X$3107 \$438 VIA_via2_5
X$3108 \$438 VIA_via2_5
X$3109 \$438 VIA_via1_4
X$3110 \$438 VIA_via1_4
X$3111 \$439 VIA_via2_5
X$3112 \$439 VIA_via2_5
X$3113 \$439 VIA_via1_4
X$3114 \$439 VIA_via1_4
X$3115 \$448 VIA_via2_5
X$3116 \$448 VIA_via1_4
X$3117 \$448 VIA_via2_5
X$3118 \$448 VIA_via1_4
X$3119 \$458 VIA_via2_5
X$3120 \$458 VIA_via1_4
X$3121 \$458 VIA_via1_4
X$3122 \$458 VIA_via2_5
X$3123 \$471 VIA_via2_5
X$3124 \$471 VIA_via2_5
X$3125 \$471 VIA_via2_5
X$3126 \$471 VIA_via2_5
X$3127 \$471 VIA_via1_4
X$3128 \$471 VIA_via1_4
X$3129 \$471 VIA_via1_4
X$3130 \$471 VIA_via2_5
X$3131 \$474 VIA_via2_5
X$3132 \$474 VIA_via2_5
X$3133 \$474 VIA_via1_4
X$3134 \$474 VIA_via2_5
X$3135 \$474 VIA_via1_4
X$3136 \$474 VIA_via1_4
X$3137 \$474 VIA_via2_5
X$3138 \$479 VIA_via2_5
X$3139 \$479 VIA_via2_5
X$3140 \$479 VIA_via1_4
X$3141 \$479 VIA_via1_4
X$3142 \$482 VIA_via2_5
X$3143 \$482 VIA_via2_5
X$3144 \$482 VIA_via1_4
X$3145 \$482 VIA_via1_4
X$3146 \$482 VIA_via1_4
X$3147 zero_flag VIA_via2_5
X$3148 zero_flag VIA_via2_5
X$3149 zero_flag VIA_via1_4
X$3150 zero_flag VIA_via2_5
X$3151 overflow_flag VIA_via2_5
X$3152 overflow_flag VIA_via2_5
X$3153 overflow_flag VIA_via1_4
X$3154 overflow_flag VIA_via2_5
X$3155 \$486 VIA_via1_4
X$3156 \$486 VIA_via2_5
X$3157 \$486 VIA_via1_4
X$3158 \$486 VIA_via2_5
X$3159 \$487 VIA_via2_5
X$3160 \$487 VIA_via1_4
X$3161 \$487 VIA_via2_5
X$3162 \$487 VIA_via1_4
X$3163 \$490 VIA_via2_5
X$3164 \$490 VIA_via1_4
X$3165 \$490 VIA_via1_4
X$3166 \$490 VIA_via2_5
X$3167 \$494 VIA_via1_4
X$3168 \$494 VIA_via2_5
X$3169 \$494 VIA_via1_4
X$3170 \$494 VIA_via2_5
X$3171 \$496 VIA_via1_4
X$3172 \$496 VIA_via2_5
X$3173 \$496 VIA_via1_4
X$3174 \$496 VIA_via2_5
X$3175 \$502 VIA_via1_4
X$3176 \$502 VIA_via2_5
X$3177 \$502 VIA_via1_4
X$3178 \$502 VIA_via2_5
X$3179 \$509 VIA_via2_5
X$3180 \$509 VIA_via1_4
X$3181 \$509 VIA_via2_5
X$3182 \$509 VIA_via1_4
X$3183 \$511 VIA_via1_4
X$3184 \$511 VIA_via2_5
X$3185 \$511 VIA_via1_4
X$3186 \$511 VIA_via2_5
X$3187 \$523 VIA_via1_4
X$3188 \$523 VIA_via2_5
X$3189 \$523 VIA_via1_4
X$3190 \$523 VIA_via2_5
X$3191 b[7] VIA_via2_5
X$3192 b[7] VIA_via1_4
X$3193 b[6] VIA_via2_5
X$3194 b[6] VIA_via1_4
X$3195 \$533 VIA_via1_4
X$3196 \$533 VIA_via2_5
X$3197 \$533 VIA_via1_4
X$3198 \$533 VIA_via1_4
X$3199 \$533 VIA_via2_5
X$3200 \$534 VIA_via1_4
X$3201 \$534 VIA_via2_5
X$3202 \$534 VIA_via1_4
X$3203 \$534 VIA_via2_5
X$3204 \$534 VIA_via1_4
X$3205 \$545 VIA_via2_5
X$3206 \$545 VIA_via2_5
X$3207 \$545 VIA_via1_4
X$3208 \$545 VIA_via1_4
X$3209 \$545 VIA_via2_5
X$3210 \$545 VIA_via1_4
X$3211 \$545 VIA_via2_5
X$3212 \$545 VIA_via1_4
X$3213 \$545 VIA_via2_5
X$3214 \$549 VIA_via2_5
X$3215 \$549 VIA_via2_5
X$3216 \$549 VIA_via2_5
X$3217 \$549 VIA_via2_5
X$3218 \$549 VIA_via2_5
X$3219 \$549 VIA_via2_5
X$3220 \$549 VIA_via2_5
X$3221 \$549 VIA_via1_4
X$3222 \$549 VIA_via2_5
X$3223 \$549 VIA_via1_4
X$3224 \$549 VIA_via1_4
X$3225 \$549 VIA_via2_5
X$3226 \$549 VIA_via1_4
X$3227 \$549 VIA_via2_5
X$3228 \$549 VIA_via1_4
X$3229 \$549 VIA_via1_4
X$3230 \$549 VIA_via1_4
X$3231 \$551 VIA_via2_5
X$3232 \$551 VIA_via2_5
X$3233 \$551 VIA_via1_4
X$3234 \$551 VIA_via2_5
X$3235 \$551 VIA_via1_4
X$3236 \$551 VIA_via1_4
X$3237 \$552 VIA_via2_5
X$3238 \$552 VIA_via2_5
X$3239 \$552 VIA_via2_5
X$3240 \$552 VIA_via2_5
X$3241 \$552 VIA_via3_2
X$3242 \$552 VIA_via2_5
X$3243 \$552 VIA_via3_2
X$3244 \$552 VIA_via2_5
X$3245 \$552 VIA_via1_4
X$3246 \$552 VIA_via1_4
X$3247 \$552 VIA_via2_5
X$3248 \$552 VIA_via1_4
X$3249 \$552 VIA_via1_4
X$3250 \$554 VIA_via2_5
X$3251 \$554 VIA_via2_5
X$3252 \$554 VIA_via2_5
X$3253 \$554 VIA_via2_5
X$3254 \$554 VIA_via2_5
X$3255 \$554 VIA_via2_5
X$3256 \$554 VIA_via1_4
X$3257 \$554 VIA_via1_4
X$3258 \$554 VIA_via2_5
X$3259 \$554 VIA_via1_4
X$3260 \$554 VIA_via1_4
X$3261 \$554 VIA_via1_4
X$3262 \$554 VIA_via1_4
X$3263 \$554 VIA_via1_4
X$3264 \$554 VIA_via2_5
X$3265 \$555 VIA_via1_4
X$3266 \$555 VIA_via1_4
X$3267 \$557 VIA_via2_5
X$3268 \$557 VIA_via1_4
X$3269 \$557 VIA_via1_4
X$3270 \$557 VIA_via2_5
X$3271 \$557 VIA_via1_4
X$3272 \$557 VIA_via2_5
X$3273 \$557 VIA_via1_4
X$3274 \$557 VIA_via1_4
X$3275 \$557 VIA_via1_4
X$3276 \$557 VIA_via1_4
X$3277 \$557 VIA_via1_4
X$3278 \$557 VIA_via1_4
X$3279 \$557 VIA_via2_5
X$3280 \$558 VIA_via2_5
X$3281 \$558 VIA_via1_4
X$3282 \$558 VIA_via2_5
X$3283 \$558 VIA_via1_4
X$3284 \$559 VIA_via2_5
X$3285 \$559 VIA_via2_5
X$3286 \$559 VIA_via1_4
X$3287 \$559 VIA_via1_4
X$3288 result[2] VIA_via2_5
X$3289 result[2] VIA_via2_5
X$3290 result[2] VIA_via2_5
X$3291 result[2] VIA_via1_4
X$3292 result[0] VIA_via2_5
X$3293 result[0] VIA_via2_5
X$3294 result[0] VIA_via1_4
X$3295 result[0] VIA_via2_5
X$3296 result[3] VIA_via2_5
X$3297 result[3] VIA_via2_5
X$3298 result[3] VIA_via1_4
X$3299 result[3] VIA_via2_5
X$3300 result[1] VIA_via2_5
X$3301 result[1] VIA_via1_4
X$3302 \$572 VIA_via2_5
X$3303 \$572 VIA_via1_4
X$3304 \$572 VIA_via2_5
X$3305 \$572 VIA_via1_4
X$3306 \$573 VIA_via2_5
X$3307 \$573 VIA_via1_4
X$3308 \$573 VIA_via2_5
X$3309 \$573 VIA_via1_4
X$3310 \$574 VIA_via2_5
X$3311 \$574 VIA_via2_5
X$3312 \$574 VIA_via2_5
X$3313 \$574 VIA_via1_4
X$3314 \$574 VIA_via2_5
X$3315 \$574 VIA_via1_4
X$3316 \$574 VIA_via2_5
X$3317 \$574 VIA_via1_4
X$3318 \$585 VIA_via2_5
X$3319 \$585 VIA_via1_4
X$3320 \$585 VIA_via2_5
X$3321 \$585 VIA_via1_4
X$3322 \$586 VIA_via2_5
X$3323 \$586 VIA_via2_5
X$3324 \$586 VIA_via1_4
X$3325 \$586 VIA_via1_4
X$3326 \$593 VIA_via2_5
X$3327 \$593 VIA_via2_5
X$3328 \$593 VIA_via2_5
X$3329 \$593 VIA_via1_4
X$3330 \$593 VIA_via2_5
X$3331 \$593 VIA_via1_4
X$3332 \$595 VIA_via2_5
X$3333 \$595 VIA_via1_4
X$3334 \$595 VIA_via1_4
X$3335 \$595 VIA_via2_5
X$3336 \$599 VIA_via2_5
X$3337 \$599 VIA_via2_5
X$3338 \$599 VIA_via1_4
X$3339 \$599 VIA_via1_4
X$3340 \$606 VIA_via3_2
X$3341 \$606 VIA_via3_2
X$3342 \$606 VIA_via2_5
X$3343 \$606 VIA_via2_5
X$3344 \$606 VIA_via2_5
X$3345 \$606 VIA_via2_5
X$3346 \$606 VIA_via2_5
X$3347 \$606 VIA_via1_4
X$3348 \$606 VIA_via1_4
X$3349 \$606 VIA_via1_4
X$3350 \$606 VIA_via1_4
X$3351 \$612 VIA_via1_4
X$3352 \$612 VIA_via1_4
X$3353 \$614 VIA_via2_5
X$3354 \$614 VIA_via2_5
X$3355 \$614 VIA_via2_5
X$3356 \$614 VIA_via1_4
X$3357 \$614 VIA_via1_4
X$3358 \$614 VIA_via1_4
X$3359 \$619 VIA_via1_4
X$3360 \$619 VIA_via1_4
X$3361 \$620 VIA_via2_5
X$3362 \$620 VIA_via1_4
X$3363 \$620 VIA_via1_4
X$3364 \$620 VIA_via2_5
X$3365 \$620 VIA_via1_4
X$3366 \$620 VIA_via2_5
X$3367 \$626 VIA_via1_4
X$3368 \$626 VIA_via1_4
X$3369 \$627 VIA_via1_4
X$3370 \$627 VIA_via1_4
X$3371 \$629 VIA_via1_4
X$3372 \$629 VIA_via1_4
X$3373 \$630 VIA_via2_5
X$3374 \$630 VIA_via1_4
X$3375 \$630 VIA_via1_4
X$3376 \$630 VIA_via2_5
X$3377 result[7] VIA_via2_5
X$3378 result[7] VIA_via1_4
X$3379 result[4] VIA_via1_4
X$3380 result[4] VIA_via2_5
X$3381 result[6] VIA_via2_5
X$3382 result[6] VIA_via2_5
X$3383 result[6] VIA_via1_4
X$3384 result[6] VIA_via2_5
X$3385 result[5] VIA_via2_5
X$3386 result[5] VIA_via2_5
X$3387 result[5] VIA_via1_4
X$3388 result[5] VIA_via2_5
X$3389 \$645 VIA_via2_5
X$3390 \$645 VIA_via2_5
X$3391 \$645 VIA_via1_4
X$3392 \$645 VIA_via1_4
X$3393 \$661 VIA_via1_4
X$3394 \$661 VIA_via1_4
X$3395 \$680 VIA_via1_4
X$3396 \$680 VIA_via2_5
X$3397 \$680 VIA_via1_4
X$3398 \$680 VIA_via2_5
X$3399 \$683 VIA_via2_5
X$3400 \$683 VIA_via1_4
X$3401 \$683 VIA_via1_4
X$3402 \$683 VIA_via2_5
X$3403 \$686 VIA_via2_5
X$3404 \$686 VIA_via2_5
X$3405 \$686 VIA_via1_4
X$3406 \$686 VIA_via1_4
X$3407 \$689 VIA_via1_4
X$3408 \$689 VIA_via2_5
X$3409 \$689 VIA_via1_4
X$3410 \$689 VIA_via2_5
X$3411 \$690 VIA_via2_5
X$3412 \$690 VIA_via1_4
X$3413 \$690 VIA_via2_5
X$3414 \$690 VIA_via1_4
X$3415 \$691 VIA_via1_4
X$3416 \$691 VIA_via2_5
X$3417 \$691 VIA_via1_4
X$3418 \$691 VIA_via2_5
X$3419 \$698 VIA_via1_4
X$3420 \$698 VIA_via2_5
X$3421 \$698 VIA_via1_4
X$3422 \$698 VIA_via2_5
X$3423 \$705 VIA_via1_4
X$3424 \$705 VIA_via2_5
X$3425 \$705 VIA_via1_4
X$3426 \$705 VIA_via2_5
X$3427 \$708 VIA_via2_5
X$3428 \$708 VIA_via1_4
X$3429 \$708 VIA_via2_5
X$3430 \$708 VIA_via1_4
X$3431 \$709 VIA_via2_5
X$3432 \$709 VIA_via1_4
X$3433 \$709 VIA_via2_5
X$3434 \$709 VIA_via1_4
X$3435 \$710 VIA_via1_4
X$3436 \$710 VIA_via2_5
X$3437 \$710 VIA_via1_4
X$3438 \$710 VIA_via2_5
X$3439 \$711 VIA_via2_5
X$3440 \$711 VIA_via1_4
X$3441 \$711 VIA_via2_5
X$3442 \$711 VIA_via1_4
X$3443 \$714 VIA_via1_4
X$3444 \$714 VIA_via2_5
X$3445 \$714 VIA_via1_4
X$3446 \$714 VIA_via2_5
X$3447 \$720 VIA_via2_5
X$3448 \$720 VIA_via1_4
X$3449 \$720 VIA_via2_5
X$3450 \$720 VIA_via1_4
X$3451 \$723 VIA_via1_4
X$3452 \$723 VIA_via2_5
X$3453 \$723 VIA_via1_4
X$3454 \$723 VIA_via2_5
X$3455 \$732 VIA_via1_4
X$3456 \$732 VIA_via2_5
X$3457 \$732 VIA_via1_4
X$3458 \$732 VIA_via2_5
X$3459 \$733 VIA_via1_4
X$3460 \$733 VIA_via2_5
X$3461 \$733 VIA_via1_4
X$3462 \$733 VIA_via2_5
X$3463 \$735 VIA_via2_5
X$3464 \$735 VIA_via1_4
X$3465 \$735 VIA_via2_5
X$3466 \$735 VIA_via1_4
X$3467 \$737 VIA_via2_5
X$3468 \$737 VIA_via2_5
X$3469 \$737 VIA_via1_4
X$3470 \$737 VIA_via1_4
X$3471 \$741 VIA_via2_5
X$3472 \$741 VIA_via1_4
X$3473 \$741 VIA_via2_5
X$3474 \$741 VIA_via1_4
X$3475 \$744 VIA_via2_5
X$3476 \$744 VIA_via1_4
X$3477 \$744 VIA_via2_5
X$3478 \$744 VIA_via1_4
X$3479 \$746 VIA_via1_4
X$3480 \$746 VIA_via2_5
X$3481 \$746 VIA_via1_4
X$3482 \$746 VIA_via2_5
X$3483 \$747 VIA_via1_4
X$3484 \$747 VIA_via2_5
X$3485 \$747 VIA_via1_4
X$3486 \$747 VIA_via2_5
X$3487 \$750 VIA_via1_7
X$3488 \$750 VIA_via1_7
X$3489 \$750 VIA_via1_4
X$3490 \$750 VIA_via1_4
X$3491 \$753 VIA_via2_5
X$3492 \$753 VIA_via2_5
X$3493 \$753 VIA_via1_4
X$3494 \$753 VIA_via1_4
X$3495 \$758 VIA_via2_5
X$3496 \$758 VIA_via1_4
X$3497 \$758 VIA_via2_5
X$3498 \$758 VIA_via1_4
X$3499 \$769 VIA_via1_4
X$3500 \$769 VIA_via2_5
X$3501 \$769 VIA_via1_4
X$3502 \$769 VIA_via2_5
X$3503 \$769 VIA_via1_4
X$3504 \$769 VIA_via1_4
X$3505 \$769 VIA_via2_5
X$3506 \$769 VIA_via1_4
X$3507 \$770 VIA_via2_5
X$3508 \$770 VIA_via2_5
X$3509 \$770 VIA_via1_4
X$3510 \$770 VIA_via1_4
X$3511 \$770 VIA_via1_4
X$3512 \$770 VIA_via1_4
X$3513 \$772 VIA_via1_4
X$3514 \$772 VIA_via2_5
X$3515 \$772 VIA_via1_4
X$3516 \$772 VIA_via1_4
X$3517 \$772 VIA_via2_5
X$3518 \$772 VIA_via1_4
X$3519 \$775 VIA_via2_5
X$3520 \$775 VIA_via2_5
X$3521 \$775 VIA_via1_4
X$3522 \$775 VIA_via1_4
X$3523 \$777 VIA_via2_5
X$3524 \$777 VIA_via1_4
X$3525 \$777 VIA_via1_4
X$3526 \$777 VIA_via2_5
X$3527 \$778 VIA_via1_4
X$3528 \$778 VIA_via1_4
X$3529 \$779 VIA_via2_5
X$3530 \$779 VIA_via1_4
X$3531 \$779 VIA_via2_5
X$3532 \$779 VIA_via1_4
X$3533 \$779 VIA_via2_5
X$3534 \$779 VIA_via1_4
X$3535 \$780 VIA_via1_4
X$3536 \$780 VIA_via2_5
X$3537 \$780 VIA_via1_4
X$3538 \$780 VIA_via2_5
X$3539 \$780 VIA_via1_4
X$3540 \$781 VIA_via1_4
X$3541 \$781 VIA_via2_5
X$3542 \$781 VIA_via1_4
X$3543 \$781 VIA_via2_5
X$3544 \$781 VIA_via1_4
X$3545 \$783 VIA_via2_5
X$3546 \$783 VIA_via1_4
X$3547 \$783 VIA_via1_4
X$3548 \$783 VIA_via2_5
X$3549 \$794 VIA_via2_5
X$3550 \$794 VIA_via1_4
X$3551 \$794 VIA_via2_5
X$3552 \$794 VIA_via1_4
X$3553 \$795 VIA_via2_5
X$3554 \$795 VIA_via2_5
X$3555 \$795 VIA_via1_4
X$3556 \$795 VIA_via1_4
X$3557 \$801 VIA_via2_5
X$3558 \$801 VIA_via2_5
X$3559 \$801 VIA_via1_4
X$3560 \$801 VIA_via1_4
X$3561 \$803 VIA_via1_7
X$3562 \$803 VIA_via2_5
X$3563 \$803 VIA_via2_5
X$3564 \$803 VIA_via1_4
X$3565 \$803 VIA_via1_4
X$3566 \$808 VIA_via2_5
X$3567 \$808 VIA_via1_4
X$3568 \$808 VIA_via1_4
X$3569 \$808 VIA_via2_5
X$3570 \$809 VIA_via2_5
X$3571 \$809 VIA_via1_4
X$3572 \$809 VIA_via1_4
X$3573 \$809 VIA_via2_5
X$3574 \$811 VIA_via2_5
X$3575 \$811 VIA_via2_5
X$3576 \$811 VIA_via1_4
X$3577 \$811 VIA_via1_4
X$3578 \$811 VIA_via1_4
X$3579 \$818 VIA_via2_5
X$3580 \$818 VIA_via2_5
X$3581 \$818 VIA_via2_5
X$3582 \$818 VIA_via1_4
X$3583 \$818 VIA_via1_4
X$3584 \$818 VIA_via2_5
X$3585 \$818 VIA_via1_4
X$3586 \$819 VIA_via2_5
X$3587 \$819 VIA_via1_4
X$3588 \$819 VIA_via1_4
X$3589 \$819 VIA_via2_5
X$3590 \$825 VIA_via2_5
X$3591 \$825 VIA_via2_5
X$3592 \$825 VIA_via2_5
X$3593 \$825 VIA_via2_5
X$3594 \$825 VIA_via2_5
X$3595 \$825 VIA_via2_5
X$3596 \$825 VIA_via2_5
X$3597 \$825 VIA_via1_4
X$3598 \$825 VIA_via1_4
X$3599 \$825 VIA_via1_4
X$3600 \$825 VIA_via2_5
X$3601 \$825 VIA_via1_4
X$3602 \$825 VIA_via1_4
X$3603 \$825 VIA_via1_4
X$3604 \$825 VIA_via1_4
X$3605 \$827 VIA_via1_7
X$3606 \$827 VIA_via2_5
X$3607 \$827 VIA_via2_5
X$3608 \$827 VIA_via1_7
X$3609 \$827 VIA_via2_5
X$3610 \$827 VIA_via1_4
X$3611 \$827 VIA_via1_4
X$3612 \$827 VIA_via1_4
X$3613 \$827 VIA_via1_4
X$3614 \$833 VIA_via2_5
X$3615 \$833 VIA_via2_5
X$3616 \$833 VIA_via1_4
X$3617 \$833 VIA_via1_4
X$3618 \$833 VIA_via1_4
X$3619 \$838 VIA_via1_4
X$3620 \$838 VIA_via1_4
X$3621 \$839 VIA_via2_5
X$3622 \$839 VIA_via1_4
X$3623 \$839 VIA_via1_4
X$3624 \$839 VIA_via1_4
X$3625 \$839 VIA_via2_5
X$3626 \$840 VIA_via1_4
X$3627 \$840 VIA_via1_4
X$3628 \$841 VIA_via2_5
X$3629 \$841 VIA_via2_5
X$3630 \$841 VIA_via1_4
X$3631 \$841 VIA_via1_4
X$3632 \$842 VIA_via1_4
X$3633 \$842 VIA_via2_5
X$3634 \$842 VIA_via1_4
X$3635 \$842 VIA_via2_5
X$3636 \$843 VIA_via1_4
X$3637 \$843 VIA_via1_4
X$3638 \$844 VIA_via1_4
X$3639 \$844 VIA_via1_4
X$3640 \$845 VIA_via2_5
X$3641 \$845 VIA_via2_5
X$3642 \$845 VIA_via1_4
X$3643 \$845 VIA_via1_4
X$3644 \$849 VIA_via1_4
X$3645 \$849 VIA_via2_5
X$3646 \$849 VIA_via1_4
X$3647 \$849 VIA_via2_5
X$3648 \$850 VIA_via2_5
X$3649 \$850 VIA_via2_5
X$3650 \$850 VIA_via1_4
X$3651 \$850 VIA_via1_4
X$3652 \$855 VIA_via2_5
X$3653 \$855 VIA_via2_5
X$3654 \$855 VIA_via1_4
X$3655 \$855 VIA_via1_4
X$3656 \$856 VIA_via2_5
X$3657 \$856 VIA_via1_4
X$3658 \$856 VIA_via2_5
X$3659 \$856 VIA_via1_4
X$3660 \$857 VIA_via2_5
X$3661 \$857 VIA_via1_4
X$3662 \$857 VIA_via2_5
X$3663 \$857 VIA_via1_4
X$3664 \$858 VIA_via2_5
X$3665 \$858 VIA_via2_5
X$3666 \$858 VIA_via1_4
X$3667 \$858 VIA_via1_4
X$3668 \$860 VIA_via2_5
X$3669 \$860 VIA_via1_4
X$3670 \$860 VIA_via1_4
X$3671 \$860 VIA_via2_5
X$3672 \$861 VIA_via2_5
X$3673 \$861 VIA_via1_4
X$3674 \$861 VIA_via2_5
X$3675 \$861 VIA_via1_4
X$3676 \$862 VIA_via1_4
X$3677 \$862 VIA_via2_5
X$3678 \$862 VIA_via1_4
X$3679 \$862 VIA_via2_5
X$3680 \$866 VIA_via2_5
X$3681 \$866 VIA_via1_4
X$3682 \$866 VIA_via2_5
X$3683 \$866 VIA_via1_4
X$3684 \$869 VIA_via2_5
X$3685 \$869 VIA_via2_5
X$3686 \$869 VIA_via2_5
X$3687 \$869 VIA_via2_5
X$3688 \$869 VIA_via1_4
X$3689 \$869 VIA_via1_4
X$3690 \$869 VIA_via1_4
X$3691 \$869 VIA_via1_4
X$3692 \$869 VIA_via2_5
X$3693 \$869 VIA_via1_4
X$3694 \$879 VIA_via1_4
X$3695 \$879 VIA_via2_5
X$3696 \$879 VIA_via1_4
X$3697 \$879 VIA_via2_5
X$3698 \$893 VIA_via2_5
X$3699 \$893 VIA_via2_5
X$3700 \$893 VIA_via2_5
X$3701 \$893 VIA_via2_5
X$3702 \$893 VIA_via2_5
X$3703 \$893 VIA_via2_5
X$3704 \$893 VIA_via2_5
X$3705 \$893 VIA_via2_5
X$3706 \$893 VIA_via2_5
X$3707 \$893 VIA_via1_4
X$3708 \$893 VIA_via1_4
X$3709 \$893 VIA_via2_5
X$3710 \$893 VIA_via1_4
X$3711 \$893 VIA_via1_4
X$3712 \$893 VIA_via1_4
X$3713 \$893 VIA_via1_4
X$3714 \$893 VIA_via1_4
X$3715 \$893 VIA_via1_4
X$3716 \$893 VIA_via1_4
X$3717 \$895 VIA_via2_5
X$3718 \$895 VIA_via2_5
X$3719 \$895 VIA_via1_4
X$3720 \$895 VIA_via2_5
X$3721 \$895 VIA_via1_4
X$3722 \$895 VIA_via2_5
X$3723 \$895 VIA_via1_4
X$3724 \$895 VIA_via1_4
X$3725 \$895 VIA_via2_5
X$3726 \$896 VIA_via2_5
X$3727 \$896 VIA_via2_5
X$3728 \$896 VIA_via1_4
X$3729 \$896 VIA_via1_4
X$3730 \$896 VIA_via1_4
X$3731 \$896 VIA_via2_5
X$3732 \$896 VIA_via1_4
X$3733 \$896 VIA_via2_5
X$3734 \$896 VIA_via1_4
X$3735 \$896 VIA_via1_4
X$3736 \$896 VIA_via2_5
X$3737 \$896 VIA_via1_4
X$3738 \$896 VIA_via2_5
X$3739 \$896 VIA_via1_4
X$3740 \$896 VIA_via1_4
X$3741 \$903 VIA_via2_5
X$3742 \$903 VIA_via1_4
X$3743 \$903 VIA_via1_4
X$3744 \$903 VIA_via2_5
X$3745 \$904 VIA_via1_4
X$3746 \$904 VIA_via1_4
X$3747 \$909 VIA_via2_5
X$3748 \$909 VIA_via2_5
X$3749 \$909 VIA_via2_5
X$3750 \$909 VIA_via2_5
X$3751 \$909 VIA_via1_4
X$3752 \$909 VIA_via1_4
X$3753 \$909 VIA_via1_4
X$3754 \$909 VIA_via1_4
X$3755 \$909 VIA_via1_4
X$3756 \$913 VIA_via2_5
X$3757 \$913 VIA_via2_5
X$3758 \$913 VIA_via1_4
X$3759 \$913 VIA_via2_5
X$3760 \$913 VIA_via1_4
X$3761 \$913 VIA_via2_5
X$3762 \$913 VIA_via1_4
X$3763 \$913 VIA_via2_5
X$3764 \$913 VIA_via1_4
X$3765 \$913 VIA_via1_4
X$3766 \$913 VIA_via1_4
X$3767 \$914 VIA_via2_5
X$3768 \$914 VIA_via1_4
X$3769 \$914 VIA_via2_5
X$3770 \$914 VIA_via1_4
X$3771 \$914 VIA_via1_4
X$3772 \$914 VIA_via2_5
X$3773 \$914 VIA_via1_4
X$3774 \$917 VIA_via1_4
X$3775 \$917 VIA_via1_4
X$3776 \$918 VIA_via1_4
X$3777 \$918 VIA_via2_5
X$3778 \$918 VIA_via1_4
X$3779 \$918 VIA_via2_5
X$3780 \$918 VIA_via1_4
X$3781 \$918 VIA_via2_5
X$3782 \$919 VIA_via2_5
X$3783 \$919 VIA_via2_5
X$3784 \$919 VIA_via2_5
X$3785 \$919 VIA_via1_4
X$3786 \$919 VIA_via1_4
X$3787 \$919 VIA_via2_5
X$3788 \$919 VIA_via1_4
X$3789 \$919 VIA_via2_5
X$3790 \$919 VIA_via1_4
X$3791 \$919 VIA_via2_5
X$3792 \$921 VIA_via1_4
X$3793 \$921 VIA_via2_5
X$3794 \$921 VIA_via1_4
X$3795 \$921 VIA_via2_5
X$3796 \$921 VIA_via1_4
X$3797 \$921 VIA_via2_5
X$3798 \$921 VIA_via1_4
X$3799 \$921 VIA_via2_5
X$3800 \$921 VIA_via1_4
X$3801 \$921 VIA_via1_4
X$3802 \$921 VIA_via2_5
X$3803 \$925 VIA_via2_5
X$3804 \$925 VIA_via1_4
X$3805 \$925 VIA_via2_5
X$3806 \$925 VIA_via1_4
X$3807 \$926 VIA_via1_4
X$3808 \$926 VIA_via1_4
X$3809 \$931 VIA_via2_5
X$3810 \$931 VIA_via1_4
X$3811 \$931 VIA_via1_4
X$3812 \$931 VIA_via2_5
X$3813 \$939 VIA_via1_4
X$3814 \$939 VIA_via2_5
X$3815 \$939 VIA_via1_4
X$3816 \$939 VIA_via2_5
X$3817 \$946 VIA_via1_4
X$3818 \$946 VIA_via2_5
X$3819 \$946 VIA_via1_4
X$3820 \$946 VIA_via2_5
X$3821 \$948 VIA_via1_4
X$3822 \$948 VIA_via2_5
X$3823 \$948 VIA_via1_4
X$3824 \$948 VIA_via2_5
X$3825 \$957 VIA_via2_5
X$3826 \$957 VIA_via1_4
X$3827 \$957 VIA_via2_5
X$3828 \$957 VIA_via1_4
X$3829 \$960 VIA_via2_5
X$3830 \$960 VIA_via1_4
X$3831 \$960 VIA_via1_4
X$3832 \$960 VIA_via2_5
X$3833 \$972 VIA_via1_7
X$3834 \$972 VIA_via2_5
X$3835 \$972 VIA_via1_4
X$3836 \$972 VIA_via2_5
X$3837 \$973 VIA_via2_5
X$3838 \$973 VIA_via2_5
X$3839 \$973 VIA_via1_4
X$3840 \$973 VIA_via1_4
X$3841 \$975 VIA_via2_5
X$3842 \$975 VIA_via1_4
X$3843 \$975 VIA_via1_4
X$3844 \$975 VIA_via2_5
X$3845 \$980 VIA_via2_5
X$3846 \$980 VIA_via1_4
X$3847 \$980 VIA_via1_4
X$3848 \$980 VIA_via2_5
X$3849 \$991 VIA_via2_5
X$3850 \$991 VIA_via1_4
X$3851 \$991 VIA_via2_5
X$3852 \$991 VIA_via1_4
X$3853 \$991 VIA_via1_4
X$3854 \$991 VIA_via2_5
X$3855 \$993 VIA_via1_4
X$3856 \$993 VIA_via1_4
X$3857 \$996 VIA_via2_5
X$3858 \$996 VIA_via2_5
X$3859 \$996 VIA_via2_5
X$3860 \$996 VIA_via1_4
X$3861 \$996 VIA_via2_5
X$3862 \$996 VIA_via1_4
X$3863 \$996 VIA_via1_4
X$3864 \$996 VIA_via2_5
X$3865 \$996 VIA_via1_4
X$3866 \$996 VIA_via2_5
X$3867 \$996 VIA_via1_4
X$3868 \$996 VIA_via1_4
X$3869 \$996 VIA_via2_5
X$3870 \$998 VIA_via2_5
X$3871 \$998 VIA_via2_5
X$3872 \$998 VIA_via2_5
X$3873 \$998 VIA_via2_5
X$3874 \$998 VIA_via2_5
X$3875 \$998 VIA_via1_4
X$3876 \$998 VIA_via2_5
X$3877 \$998 VIA_via1_4
X$3878 \$998 VIA_via2_5
X$3879 \$998 VIA_via1_4
X$3880 \$998 VIA_via1_4
X$3881 \$998 VIA_via2_5
X$3882 \$998 VIA_via1_4
X$3883 \$999 VIA_via1_4
X$3884 \$999 VIA_via1_4
X$3885 \$999 VIA_via2_5
X$3886 \$999 VIA_via1_4
X$3887 \$999 VIA_via2_5
X$3888 \$999 VIA_via1_4
X$3889 \$999 VIA_via2_5
X$3890 \$999 VIA_via1_4
X$3891 \$999 VIA_via1_4
X$3892 \$1001 VIA_via1_4
X$3893 \$1001 VIA_via1_4
X$3894 \$1002 VIA_via1_4
X$3895 \$1002 VIA_via1_4
X$3896 \$1003 VIA_via2_5
X$3897 \$1003 VIA_via1_4
X$3898 \$1003 VIA_via2_5
X$3899 \$1003 VIA_via1_4
X$3900 \$1003 VIA_via2_5
X$3901 \$1003 VIA_via1_4
X$3902 \$1004 VIA_via2_5
X$3903 \$1004 VIA_via1_4
X$3904 \$1004 VIA_via2_5
X$3905 \$1004 VIA_via1_4
X$3906 \$1004 VIA_via2_5
X$3907 \$1004 VIA_via1_4
X$3908 \$1006 VIA_via2_5
X$3909 \$1006 VIA_via2_5
X$3910 \$1006 VIA_via2_5
X$3911 \$1006 VIA_via1_4
X$3912 \$1006 VIA_via1_4
X$3913 \$1006 VIA_via1_4
X$3914 \$1008 VIA_via2_5
X$3915 \$1008 VIA_via1_4
X$3916 \$1008 VIA_via1_4
X$3917 \$1008 VIA_via2_5
X$3918 \$1012 VIA_via1_4
X$3919 \$1012 VIA_via2_5
X$3920 \$1012 VIA_via1_4
X$3921 \$1012 VIA_via2_5
X$3922 \$1015 VIA_via1_4
X$3923 \$1015 VIA_via2_5
X$3924 \$1015 VIA_via1_4
X$3925 \$1015 VIA_via2_5
X$3926 \$1016 VIA_via1_4
X$3927 \$1016 VIA_via2_5
X$3928 \$1016 VIA_via1_4
X$3929 \$1016 VIA_via2_5
X$3930 \$1019 VIA_via2_5
X$3931 \$1019 VIA_via2_5
X$3932 \$1019 VIA_via1_4
X$3933 \$1019 VIA_via1_4
X$3934 clk VIA_via5_0
X$3935 clk VIA_via4_0
X$3936 clk VIA_via4_0
X$3937 clk VIA_via5_0
X$3938 clk VIA_via3_2
X$3939 clk VIA_via1_4
X$3940 clk VIA_via2_5
X$3941 \$1042 VIA_via2_5
X$3942 \$1042 VIA_via1_4
X$3943 \$1042 VIA_via2_5
X$3944 \$1042 VIA_via1_4
X$3945 \$1046 VIA_via1_4
X$3946 \$1046 VIA_via2_5
X$3947 \$1046 VIA_via1_4
X$3948 \$1046 VIA_via2_5
X$3949 \$1050 VIA_via1_7
X$3950 \$1050 VIA_via1_7
X$3951 \$1050 VIA_via2_5
X$3952 \$1050 VIA_via2_5
X$3953 \$1050 VIA_via1_4
X$3954 \$1050 VIA_via1_4
X$3955 \$1050 VIA_via1_4
X$3956 \$1050 VIA_via1_4
X$3957 \$1050 VIA_via2_5
X$3958 \$1050 VIA_via1_4
X$3959 \$1055 VIA_via2_5
X$3960 \$1055 VIA_via1_4
X$3961 \$1055 VIA_via1_4
X$3962 \$1055 VIA_via2_5
X$3963 \$1056 VIA_via2_5
X$3964 \$1056 VIA_via1_4
X$3965 \$1056 VIA_via2_5
X$3966 \$1056 VIA_via1_4
X$3967 \$1059 VIA_via1_4
X$3968 \$1059 VIA_via1_4
X$3969 \$1061 VIA_via2_5
X$3970 \$1061 VIA_via2_5
X$3971 \$1061 VIA_via1_4
X$3972 \$1061 VIA_via1_4
X$3973 \$1062 VIA_via2_5
X$3974 \$1062 VIA_via2_5
X$3975 \$1062 VIA_via1_4
X$3976 \$1062 VIA_via1_4
X$3977 \$1067 VIA_via2_5
X$3978 \$1067 VIA_via1_4
X$3979 \$1067 VIA_via2_5
X$3980 \$1067 VIA_via1_4
X$3981 \$1070 VIA_via2_5
X$3982 \$1070 VIA_via1_4
X$3983 \$1070 VIA_via1_4
X$3984 \$1070 VIA_via2_5
X$3985 \$1076 VIA_via2_5
X$3986 \$1076 VIA_via1_4
X$3987 \$1076 VIA_via2_5
X$3988 \$1076 VIA_via1_4
X$3989 \$1077 VIA_via2_5
X$3990 \$1077 VIA_via1_4
X$3991 \$1077 VIA_via2_5
X$3992 \$1077 VIA_via1_4
X$3993 \$1078 VIA_via2_5
X$3994 \$1078 VIA_via1_4
X$3995 \$1078 VIA_via1_4
X$3996 \$1078 VIA_via2_5
X$3997 \$1084 VIA_via1_4
X$3998 \$1084 VIA_via2_5
X$3999 \$1084 VIA_via1_4
X$4000 \$1084 VIA_via2_5
X$4001 \$1088 VIA_via1_4
X$4002 \$1088 VIA_via1_4
X$4003 \$1089 VIA_via2_5
X$4004 \$1089 VIA_via2_5
X$4005 \$1089 VIA_via1_4
X$4006 \$1089 VIA_via1_4
X$4007 \$1093 VIA_via2_5
X$4008 \$1093 VIA_via1_4
X$4009 \$1093 VIA_via1_4
X$4010 \$1093 VIA_via2_5
X$4011 \$1093 VIA_via1_4
X$4012 \$1093 VIA_via2_5
X$4013 \$1093 VIA_via1_4
X$4014 \$1093 VIA_via2_5
X$4015 \$1096 VIA_via2_5
X$4016 \$1096 VIA_via2_5
X$4017 \$1096 VIA_via1_4
X$4018 \$1096 VIA_via2_5
X$4019 \$1096 VIA_via1_4
X$4020 \$1096 VIA_via1_4
X$4021 \$1097 VIA_via2_5
X$4022 \$1097 VIA_via2_5
X$4023 \$1097 VIA_via1_4
X$4024 \$1097 VIA_via1_4
X$4025 \$1097 VIA_via2_5
X$4026 \$1097 VIA_via1_4
X$4027 \$1097 VIA_via1_4
X$4028 \$1097 VIA_via1_4
X$4029 \$1097 VIA_via1_4
X$4030 \$1097 VIA_via2_5
X$4031 \$1098 VIA_via1_4
X$4032 \$1098 VIA_via1_4
X$4033 \$1101 VIA_via2_5
X$4034 \$1101 VIA_via1_4
X$4035 \$1101 VIA_via2_5
X$4036 \$1101 VIA_via1_4
X$4037 \$1101 VIA_via1_4
X$4038 \$1101 VIA_via2_5
X$4039 \$1108 VIA_via4_0
X$4040 \$1108 VIA_via3_2
X$4041 \$1108 VIA_via3_2
X$4042 \$1108 VIA_via4_0
X$4043 \$1108 VIA_via3_2
X$4044 \$1108 VIA_via2_5
X$4045 \$1108 VIA_via2_5
X$4046 \$1108 VIA_via2_5
X$4047 \$1108 VIA_via2_5
X$4048 \$1108 VIA_via2_5
X$4049 \$1108 VIA_via1_4
X$4050 \$1108 VIA_via1_4
X$4051 \$1108 VIA_via2_5
X$4052 \$1108 VIA_via1_4
X$4053 \$1108 VIA_via1_4
X$4054 \$1109 VIA_via1_4
X$4055 \$1109 VIA_via1_4
X$4056 \$1111 VIA_via2_5
X$4057 \$1111 VIA_via2_5
X$4058 \$1111 VIA_via2_5
X$4059 \$1111 VIA_via1_4
X$4060 \$1111 VIA_via1_4
X$4061 \$1111 VIA_via1_4
X$4062 \$1111 VIA_via2_5
X$4063 \$1112 VIA_via1_4
X$4064 \$1112 VIA_via1_4
X$4065 \$1113 VIA_via2_5
X$4066 \$1113 VIA_via1_4
X$4067 \$1113 VIA_via2_5
X$4068 \$1113 VIA_via1_4
X$4069 \$1113 VIA_via2_5
X$4070 \$1113 VIA_via1_4
X$4071 \$1114 VIA_via1_4
X$4072 \$1114 VIA_via1_4
X$4073 \$1115 VIA_via2_5
X$4074 \$1115 VIA_via1_4
X$4075 \$1115 VIA_via1_4
X$4076 \$1115 VIA_via2_5
X$4077 \$1115 VIA_via1_4
X$4078 \$1115 VIA_via2_5
X$4079 \$1116 VIA_via2_5
X$4080 \$1116 VIA_via2_5
X$4081 \$1116 VIA_via2_5
X$4082 \$1116 VIA_via1_4
X$4083 \$1116 VIA_via1_4
X$4084 \$1116 VIA_via2_5
X$4085 \$1116 VIA_via1_4
X$4086 \$1116 VIA_via2_5
X$4087 \$1116 VIA_via1_4
X$4088 \$1116 VIA_via2_5
X$4089 \$1116 VIA_via1_4
X$4090 \$1116 VIA_via1_4
X$4091 \$1121 VIA_via1_4
X$4092 \$1121 VIA_via2_5
X$4093 \$1121 VIA_via1_4
X$4094 \$1121 VIA_via2_5
X$4095 \$1123 VIA_via1_4
X$4096 \$1123 VIA_via2_5
X$4097 \$1123 VIA_via1_4
X$4098 \$1123 VIA_via2_5
X$4099 \$1127 VIA_via1_4
X$4100 \$1127 VIA_via1_4
X$4101 \$1127 VIA_via2_5
X$4102 \$1127 VIA_via1_4
X$4103 \$1127 VIA_via2_5
X$4104 \$1137 VIA_via1_7
X$4105 \$1137 VIA_via1_7
X$4106 \$1137 VIA_via2_5
X$4107 \$1137 VIA_via2_5
X$4108 \$1137 VIA_via2_5
X$4109 \$1137 VIA_via2_5
X$4110 \$1137 VIA_via1_4
X$4111 \$1137 VIA_via1_4
X$4112 \$1137 VIA_via1_4
X$4113 \$1142 VIA_via2_5
X$4114 \$1142 VIA_via1_4
X$4115 \$1142 VIA_via1_4
X$4116 \$1142 VIA_via2_5
X$4117 rst_n VIA_via3_2
X$4118 rst_n VIA_via1_4
X$4119 rst_n VIA_via2_5
X$4120 \$1151 VIA_via1_4
X$4121 \$1151 VIA_via2_5
X$4122 \$1151 VIA_via1_4
X$4123 \$1151 VIA_via2_5
X$4124 \$1153 VIA_via2_5
X$4125 \$1153 VIA_via1_4
X$4126 \$1153 VIA_via2_5
X$4127 \$1153 VIA_via1_4
X$4128 \$1157 VIA_via1_4
X$4129 \$1157 VIA_via2_5
X$4130 \$1157 VIA_via1_4
X$4131 \$1157 VIA_via2_5
X$4132 \$1162 VIA_via2_5
X$4133 \$1162 VIA_via2_5
X$4134 \$1162 VIA_via1_4
X$4135 \$1162 VIA_via1_4
X$4136 \$1162 VIA_via2_5
X$4137 \$1162 VIA_via1_4
X$4138 \$1162 VIA_via2_5
X$4139 \$1162 VIA_via1_4
X$4140 \$1162 VIA_via2_5
X$4141 \$1171 VIA_via1_7
X$4142 \$1171 VIA_via1_7
X$4143 \$1171 VIA_via1_4
X$4144 \$1171 VIA_via1_4
X$4145 \$1177 VIA_via2_5
X$4146 \$1177 VIA_via2_5
X$4147 \$1177 VIA_via2_5
X$4148 \$1177 VIA_via1_4
X$4149 \$1177 VIA_via1_4
X$4150 \$1177 VIA_via1_4
X$4151 \$1178 VIA_via1_4
X$4152 \$1178 VIA_via1_4
X$4153 \$1182 VIA_via1_7
X$4154 \$1182 VIA_via2_5
X$4155 \$1182 VIA_via2_5
X$4156 \$1182 VIA_via2_5
X$4157 \$1182 VIA_via2_5
X$4158 \$1182 VIA_via2_5
X$4159 \$1182 VIA_via1_4
X$4160 \$1182 VIA_via1_4
X$4161 \$1182 VIA_via1_4
X$4162 \$1182 VIA_via1_4
X$4163 \$1184 VIA_via1_4
X$4164 \$1184 VIA_via2_5
X$4165 \$1184 VIA_via1_4
X$4166 \$1184 VIA_via2_5
X$4167 \$1185 VIA_via1_4
X$4168 \$1185 VIA_via1_4
X$4169 \$1186 VIA_via1_4
X$4170 \$1186 VIA_via1_4
X$4171 \$1187 VIA_via1_4
X$4172 \$1187 VIA_via1_4
X$4173 \$1188 VIA_via2_5
X$4174 \$1188 VIA_via1_4
X$4175 \$1188 VIA_via2_5
X$4176 \$1188 VIA_via1_4
X$4177 \$1193 VIA_via2_5
X$4178 \$1193 VIA_via1_4
X$4179 \$1193 VIA_via1_4
X$4180 \$1193 VIA_via2_5
X$4181 \$1195 VIA_via1_4
X$4182 \$1195 VIA_via2_5
X$4183 \$1195 VIA_via1_4
X$4184 \$1195 VIA_via2_5
X$4185 \$1208 VIA_via1_4
X$4186 \$1208 VIA_via2_5
X$4187 \$1208 VIA_via1_4
X$4188 \$1208 VIA_via2_5
X$4189 \$1217 VIA_via2_5
X$4190 \$1217 VIA_via2_5
X$4191 \$1217 VIA_via1_4
X$4192 \$1217 VIA_via2_5
X$4193 \$1217 VIA_via1_4
X$4194 \$1217 VIA_via2_5
X$4195 \$1220 VIA_via2_5
X$4196 \$1220 VIA_via1_4
X$4197 \$1220 VIA_via1_4
X$4198 \$1220 VIA_via2_5
X$4199 \$1222 VIA_via2_5
X$4200 \$1222 VIA_via2_5
X$4201 \$1222 VIA_via2_5
X$4202 \$1222 VIA_via2_5
X$4203 \$1222 VIA_via1_4
X$4204 \$1222 VIA_via1_4
X$4205 \$1222 VIA_via1_4
X$4206 \$1222 VIA_via2_5
X$4207 \$1225 VIA_via2_5
X$4208 \$1225 VIA_via1_4
X$4209 \$1225 VIA_via1_4
X$4210 \$1225 VIA_via2_5
X$4211 \$1230 VIA_via2_5
X$4212 \$1230 VIA_via1_4
X$4213 \$1230 VIA_via2_5
X$4214 \$1230 VIA_via1_4
X$4215 \$1242 VIA_via2_5
X$4216 \$1242 VIA_via1_4
X$4217 \$1242 VIA_via2_5
X$4218 \$1242 VIA_via1_4
X$4219 \$1246 VIA_via1_4
X$4220 \$1246 VIA_via1_4
X$4221 \$1253 VIA_via1_4
X$4222 \$1253 VIA_via1_4
X$4223 \$1253 VIA_via1_4
X$4224 \$1254 VIA_via2_5
X$4225 \$1254 VIA_via2_5
X$4226 \$1254 VIA_via2_5
X$4227 \$1254 VIA_via2_5
X$4228 \$1254 VIA_via2_5
X$4229 \$1254 VIA_via2_5
X$4230 \$1254 VIA_via2_5
X$4231 \$1254 VIA_via1_4
X$4232 \$1254 VIA_via2_5
X$4233 \$1254 VIA_via1_4
X$4234 \$1254 VIA_via2_5
X$4235 \$1254 VIA_via1_4
X$4236 \$1254 VIA_via1_4
X$4237 \$1254 VIA_via1_4
X$4238 \$1254 VIA_via1_4
X$4239 \$1254 VIA_via1_4
X$4240 \$1254 VIA_via1_4
X$4241 opcode[1] VIA_via3_2
X$4242 opcode[1] VIA_via2_5
X$4243 opcode[1] VIA_via2_5
X$4244 opcode[1] VIA_via2_5
X$4245 opcode[1] VIA_via1_4
X$4246 opcode[1] VIA_via2_5
X$4247 opcode[1] VIA_via1_4
X$4248 opcode[1] VIA_via1_4
X$4249 opcode[1] VIA_via1_4
X$4250 opcode[1] VIA_via2_5
X$4251 opcode[1] VIA_via1_4
X$4252 opcode[1] VIA_via1_4
X$4253 opcode[1] VIA_via2_5
X$4254 \$1258 VIA_via2_5
X$4255 \$1258 VIA_via1_4
X$4256 \$1258 VIA_via2_5
X$4257 \$1258 VIA_via1_4
X$4258 \$1258 VIA_via1_4
X$4259 \$1258 VIA_via1_4
X$4260 \$1258 VIA_via2_5
X$4261 \$1258 VIA_via1_4
X$4262 \$1258 VIA_via2_5
X$4263 \$1258 VIA_via1_4
X$4264 \$1258 VIA_via2_5
X$4265 \$1261 VIA_via2_5
X$4266 \$1261 VIA_via2_5
X$4267 \$1261 VIA_via2_5
X$4268 \$1261 VIA_via1_4
X$4269 \$1261 VIA_via2_5
X$4270 \$1261 VIA_via1_4
X$4271 \$1261 VIA_via2_5
X$4272 \$1261 VIA_via1_4
X$4273 \$1261 VIA_via1_4
X$4274 \$1265 VIA_via2_5
X$4275 \$1265 VIA_via1_4
X$4276 \$1265 VIA_via1_4
X$4277 \$1265 VIA_via2_5
X$4278 \$1270 VIA_via2_5
X$4279 \$1270 VIA_via2_5
X$4280 \$1270 VIA_via1_4
X$4281 \$1270 VIA_via1_4
X$4282 \$1279 VIA_via2_5
X$4283 \$1279 VIA_via1_4
X$4284 \$1279 VIA_via1_4
X$4285 \$1279 VIA_via2_5
X$4286 \$1283 VIA_via1_4
X$4287 \$1283 VIA_via2_5
X$4288 \$1283 VIA_via1_4
X$4289 \$1283 VIA_via2_5
X$4290 \$1291 VIA_via1_4
X$4291 \$1291 VIA_via2_5
X$4292 \$1291 VIA_via1_4
X$4293 \$1291 VIA_via2_5
X$4294 \$1298 VIA_via1_4
X$4295 \$1298 VIA_via2_5
X$4296 \$1298 VIA_via1_4
X$4297 \$1298 VIA_via2_5
X$4298 \$1305 VIA_via2_5
X$4299 \$1305 VIA_via1_4
X$4300 \$1305 VIA_via2_5
X$4301 \$1305 VIA_via1_4
X$4302 \$1314 VIA_via2_5
X$4303 \$1314 VIA_via2_5
X$4304 \$1314 VIA_via1_4
X$4305 \$1314 VIA_via2_5
X$4306 \$1314 VIA_via1_4
X$4307 \$1314 VIA_via1_4
X$4308 \$1315 VIA_via1_4
X$4309 \$1315 VIA_via1_4
X$4310 opcode[3] VIA_via3_2
X$4311 opcode[3] VIA_via2_5
X$4312 opcode[3] VIA_via2_5
X$4313 opcode[3] VIA_via1_4
X$4314 opcode[3] VIA_via2_5
X$4315 opcode[3] VIA_via1_4
X$4316 opcode[0] VIA_via3_2
X$4317 opcode[0] VIA_via1_4
X$4318 opcode[0] VIA_via2_5
X$4319 opcode[0] VIA_via1_4
X$4320 opcode[0] VIA_via2_5
X$4321 \$1319 VIA_via1_4
X$4322 \$1319 VIA_via1_4
X$4323 \$1320 VIA_via1_4
X$4324 \$1320 VIA_via1_4
X$4325 \$1338 VIA_via2_5
X$4326 \$1338 VIA_via1_4
X$4327 \$1338 VIA_via2_5
X$4328 \$1338 VIA_via1_4
X$4329 \$1339 VIA_via1_4
X$4330 \$1339 VIA_via2_5
X$4331 \$1339 VIA_via1_4
X$4332 \$1339 VIA_via2_5
X$4333 opcode[2] VIA_via3_2
X$4334 opcode[2] VIA_via1_4
X$4335 opcode[2] VIA_via2_5
.ENDS alu

.SUBCKT XNOR2_X2 A B VSS NWELL|VDD ZN PWELL
M$1 ZN A \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U
+ PD=0.77U
M$2 \$11 A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$3 NWELL|VDD B \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 \$8 B NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 ZN \$1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$6 NWELL|VDD \$1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 \$1 B NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 NWELL|VDD A \$1 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 \$6 A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$10 ZN A \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$11 \$6 B ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$12 ZN B \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
M$13 \$6 \$1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$14 VSS \$1 \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 \$12 B VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 \$1 A \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS XNOR2_X2

.SUBCKT OAI211_X2 A B C2 C1 ZN VSS NWELL|VDD PWELL
M$1 ZN A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD B ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN B NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P
+ PS=0.77U PD=0.775U
M$4 NWELL|VDD A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0441P
+ PS=0.775U PD=0.77U
M$5 \$12 C2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 ZN C1 \$12 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 \$11 C1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 NWELL|VDD C2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 \$14 A \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$10 VSS B \$14 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 \$13 B VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P
+ PS=0.555U PD=0.56U
M$12 \$5 A \$13 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.02905P
+ PS=0.56U PD=0.555U
M$13 ZN C2 \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$14 \$5 C1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN C1 \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 \$5 C2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OAI211_X2

.SUBCKT AOI21_X4 VSS ZN A B2 B1 NWELL|VDD PWELL
M$1 NWELL|VDD A \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$11 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD A \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 \$11 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 ZN B2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 \$11 B1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 ZN B1 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 \$11 B2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$9 ZN B2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$10 \$11 B1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$11 ZN B1 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$12 \$11 B2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$13 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$14 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$15 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$16 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$17 \$8 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$18 ZN B1 \$8 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$19 \$9 B1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$20 VSS B2 \$9 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$21 \$6 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$22 ZN B1 \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$23 \$7 B1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$24 VSS B2 \$7 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AOI21_X4

.SUBCKT AND3_X1 A1 A2 A3 NWELL|VDD VSS ZN PWELL
M$1 NWELL|VDD A1 \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.84U PD=0.455U
M$2 \$4 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P
+ AD=0.02205P PS=0.455U PD=0.455U
M$3 \$4 A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.77U PD=0.455U
M$4 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P
+ AD=0.06615P PS=0.77U PD=1.47U
M$5 \$10 A1 \$4 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$6 \$11 A2 \$10 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$7 VSS A3 \$11 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
M$8 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AND3_X1

.SUBCKT OR2_X2 A1 A2 VSS NWELL|VDD ZN PWELL
M$1 \$9 A1 \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A2 \$9 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD \$4 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 \$4 A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$6 VSS A2 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$7 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 VSS \$4 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OR2_X2

.SUBCKT OR2_X1 A1 A2 VSS NWELL|VDD ZN PWELL
M$1 \$9 A1 \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P
+ PS=0.84U PD=0.455U
M$2 \$9 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.77U PD=0.455U
M$3 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P
+ AD=0.06615P PS=0.77U PD=1.47U
M$4 \$4 A1 VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$5 VSS A2 \$4 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
M$6 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OR2_X1

.SUBCKT AOI221_X2 B1 B2 A C2 C1 ZN NWELL|VDD VSS PWELL
M$1 \$7 A \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD B1 \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$7 B2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD B2 \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 \$7 B1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 \$10 A \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.04725P
+ PS=0.77U PD=0.78U
M$7 ZN C2 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.04725P AD=0.0441P
+ PS=0.78U PD=0.77U
M$8 \$10 C1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$9 ZN C1 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$10 \$10 C2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$11 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$12 \$16 B1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$13 VSS B2 \$16 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$14 \$15 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN B1 \$15 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.031125P
+ PS=0.555U PD=0.565U
M$17 \$14 C2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.031125P AD=0.02905P
+ PS=0.565U PD=0.555U
M$18 ZN C1 \$14 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$19 \$13 C1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$20 VSS C2 \$13 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AOI221_X2

.SUBCKT OR3_X2 A1 A2 A3 VSS NWELL|VDD ZN PWELL
M$1 \$11 A1 \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$10 A2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD A3 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 NWELL|VDD \$4 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$6 VSS A1 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$7 \$4 A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 VSS A3 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$9 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$10 VSS \$4 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OR3_X2

.SUBCKT NAND2_X2 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 \$9 A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$6 ZN A1 \$9 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$7 \$8 A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$8 VSS A2 \$8 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NAND2_X2

.SUBCKT INV_X2 A VSS NWELL|VDD ZN PWELL
M$1 ZN A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$3 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$4 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS INV_X2

.SUBCKT OAI21_X2 A B2 B1 NWELL|VDD VSS ZN PWELL
M$1 ZN A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$10 B2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 ZN B1 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 \$11 B1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 NWELL|VDD B2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$7 VSS A \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$8 \$4 A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$9 ZN B2 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$10 \$4 B1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 ZN B1 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 \$4 B2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OAI21_X2

.SUBCKT AOI21_X2 A B2 B1 VSS ZN NWELL|VDD PWELL
M$1 NWELL|VDD A \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$5 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN B2 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$4 \$5 B1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$5 ZN B1 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$6 \$5 B2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$7 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$8 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$9 \$11 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$10 ZN B1 \$11 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 \$10 B1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 VSS B2 \$10 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AOI21_X2

.SUBCKT OR4_X1 A1 A2 A3 A4 VSS NWELL|VDD ZN PWELL
M$1 \$12 A1 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P
+ PS=0.84U PD=0.455U
M$2 \$11 A2 \$12 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P
+ PS=0.455U PD=0.455U
M$3 \$13 A3 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P
+ PS=0.455U PD=0.455U
M$4 \$13 A4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.77U PD=0.455U
M$5 ZN \$6 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P
+ AD=0.06615P PS=0.77U PD=1.47U
M$6 \$6 A1 VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$7 VSS A2 \$6 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$8 \$6 A3 VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$9 VSS A4 \$6 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
M$10 ZN \$6 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OR4_X1

.SUBCKT NAND3_X4 A2 A1 A3 VSS ZN NWELL|VDD PWELL
M$1 ZN A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 NWELL|VDD A3 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 ZN A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 NWELL|VDD A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$9 ZN A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$10 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$11 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$12 NWELL|VDD A3 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$13 \$15 A3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$14 \$14 A2 \$15 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN A1 \$14 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 \$12 A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$17 \$10 A2 \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$18 VSS A3 \$10 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$19 \$11 A3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$20 \$9 A2 \$11 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$21 ZN A1 \$9 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$22 \$16 A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$23 \$13 A2 \$16 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$24 VSS A3 \$13 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NAND3_X4

.SUBCKT NOR3_X4 VSS A1 A2 A3 ZN NWELL|VDD PWELL
M$1 ZN A1 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$8 A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$3 ZN A1 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$4 \$8 A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$5 \$6 A2 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 \$8 A2 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 \$6 A2 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 \$8 A2 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 \$6 A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$10 NWELL|VDD A3 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$11 \$6 A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$12 NWELL|VDD A3 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$13 ZN A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$14 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$17 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$18 VSS A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$19 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$20 VSS A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
M$21 ZN A3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$22 VSS A3 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$23 ZN A3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$24 VSS A3 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NOR3_X4

.SUBCKT OR2_X4 A2 A1 VSS ZN NWELL|VDD PWELL
M$1 \$10 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$4 A1 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$9 A1 \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A2 \$9 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 NWELL|VDD \$4 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 NWELL|VDD \$4 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 \$4 A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$10 VSS A1 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 \$4 A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 VSS A2 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$13 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$14 VSS \$4 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 VSS \$4 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OR2_X4

.SUBCKT NAND2_X4 A2 A1 VSS ZN NWELL|VDD PWELL
M$1 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 ZN A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$7 ZN A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$8 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 VSS A2 \$3 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$10 \$3 A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 VSS A2 \$3 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 \$3 A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$13 ZN A1 \$3 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$14 \$3 A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN A1 \$3 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 \$3 A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NAND2_X4

.SUBCKT NOR4_X1 A4 A3 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 \$12 A4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$11 A3 \$12 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$10 A2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 ZN A1 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 ZN A4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$6 VSS A3 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$7 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$8 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NOR4_X1

.SUBCKT NAND4_X1 A4 A3 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 ZN A4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A3 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 \$12 A4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$6 \$11 A3 \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$7 \$10 A2 \$11 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 ZN A1 \$10 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NAND4_X1

.SUBCKT CLKBUF_X3 A VSS NWELL|VDD Z PWELL
M$1 NWELL|VDD A \$2 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD \$2 Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 VSS A \$2 PWELL NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U
+ PD=0.335U
M$6 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.01365P PS=0.335U
+ PD=0.335U
M$7 VSS \$2 Z PWELL NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.01365P PS=0.335U
+ PD=0.335U
M$8 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.020475P
+ PS=0.335U PD=0.6U
.ENDS CLKBUF_X3

.SUBCKT CLKBUF_X1 A VSS NWELL|VDD Z PWELL
M$1 \$2 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.033075P PS=0.77U PD=0.84U
M$2 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P
+ PS=0.77U PD=1.47U
M$3 VSS A \$2 PWELL NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U
+ PD=0.335U
M$4 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P
+ PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

.SUBCKT BUF_X4 A NWELL|VDD Z VSS PWELL
M$1 \$2 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A \$2 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD \$2 Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 NWELL|VDD \$2 Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$7 \$2 A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$8 VSS A \$2 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$9 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$10 VSS \$2 Z PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 VSS \$2 Z PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS BUF_X4

.SUBCKT BUF_X1 A VSS NWELL|VDD Z PWELL
M$1 \$2 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.033075P PS=0.77U PD=0.84U
M$2 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P
+ PS=0.77U PD=1.47U
M$3 VSS A \$2 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U
+ PD=0.555U
M$4 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS BUF_X1

.SUBCKT CLKBUF_X2 A VSS NWELL|VDD Z PWELL
M$1 NWELL|VDD A \$2 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD \$2 Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$4 VSS A \$2 PWELL NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U
+ PD=0.335U
M$5 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.01365P PS=0.335U
+ PD=0.335U
M$6 VSS \$2 Z PWELL NMOS_VTL L=0.05U W=0.195U AS=0.01365P AD=0.020475P
+ PS=0.335U PD=0.6U
.ENDS CLKBUF_X2

.SUBCKT BUF_X2 A VSS NWELL|VDD Z PWELL
M$1 NWELL|VDD A \$2 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 Z \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD \$2 Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$4 VSS A \$2 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$5 Z \$2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$6 VSS \$2 Z PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS BUF_X2

.SUBCKT DFF_X2 VSS D CK Q NWELL|VDD PWELL
M$1 QN \$9 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD \$9 QN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 Q \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD \$2 Q NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 NWELL|VDD \$7 \$3 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.014175P PS=0.84U PD=0.455U
M$6 \$18 \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.09U AS=0.014175P
+ AD=0.0063P PS=0.455U PD=0.23U
M$7 \$18 \$7 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P
+ PS=0.56U PD=0.23U
M$8 \$19 \$3 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.42U AS=0.01785P AD=0.0294P
+ PS=0.56U PD=0.56U
M$9 NWELL|VDD D \$19 NWELL|VDD PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P
+ PS=0.56U PD=0.56U
M$10 \$4 \$5 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.025725P
+ AD=0.0567P PS=0.56U PD=0.99U
M$11 \$21 \$3 \$9 NWELL|VDD PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P
+ PS=0.455U PD=0.23U
M$12 \$21 \$2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.09U AS=0.0252P
+ AD=0.0063P PS=0.77U PD=0.23U
M$13 NWELL|VDD CK \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.84U PD=0.455U
M$14 \$20 \$5 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P
+ AD=0.02205P PS=0.455U PD=0.455U
M$15 \$9 \$7 \$20 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P
+ PS=0.455U PD=0.455U
M$16 \$2 \$9 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0252P
+ AD=0.06615P PS=0.77U PD=1.47U
M$17 QN \$9 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$18 VSS \$9 QN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$19 Q \$2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$20 VSS \$2 Q PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
M$21 \$13 \$4 VSS PWELL NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U
+ PD=0.23U
M$22 \$13 \$3 \$5 PWELL NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P
+ PS=0.415U PD=0.23U
M$23 \$4 \$5 VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P
+ PS=0.415U PD=0.63U
M$24 \$14 \$7 \$5 PWELL NMOS_VTL L=0.05U W=0.275U AS=0.012775P AD=0.01925P
+ PS=0.415U PD=0.415U
M$25 VSS D \$14 PWELL NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P
+ PS=0.415U PD=0.415U
M$26 VSS \$7 \$3 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U
+ PD=0.35U
M$27 VSS CK \$7 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$28 \$15 \$5 VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$29 \$9 \$3 \$15 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U
+ PD=0.35U
M$30 \$16 \$7 \$9 PWELL NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U
+ PD=0.23U
M$31 \$16 \$2 VSS PWELL NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P
+ PS=0.555U PD=0.23U
M$32 \$2 \$9 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS DFF_X2

.SUBCKT OAI22_X1 B2 B1 A1 A2 NWELL|VDD VSS ZN PWELL
M$1 \$12 B2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN B1 \$12 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$11 A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 VSS B2 \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$6 \$5 B1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$7 ZN A1 \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$8 \$5 A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OAI22_X1

.SUBCKT OAI221_X1 B2 B1 A C2 C1 NWELL|VDD VSS ZN PWELL
M$1 \$14 B2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN B1 \$14 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 \$13 C2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 ZN C1 \$13 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$6 VSS B2 \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$7 \$6 B1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 \$10 A \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$9 ZN C2 \$10 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$10 \$10 C1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OAI221_X1

.SUBCKT AOI22_X1 B2 B1 A1 A2 VSS NWELL|VDD ZN PWELL
M$1 NWELL|VDD B2 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$6 B1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A1 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$4 \$6 A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 \$12 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$6 ZN B1 \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$7 \$11 A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 VSS A2 \$11 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AOI22_X1

.SUBCKT AOI221_X1 B2 B1 A C2 C1 VSS NWELL|VDD ZN PWELL
M$1 NWELL|VDD B2 \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$7 B1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$10 A \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 ZN C2 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 \$10 C1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$6 \$14 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$7 ZN B1 \$14 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$9 \$13 C2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$10 ZN C1 \$13 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AOI221_X1

.SUBCKT AOI21_X1 A B2 B1 VSS ZN NWELL|VDD PWELL
M$1 ZN B2 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$5 B1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$3 NWELL|VDD A \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$4 \$10 B2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$5 ZN B1 \$10 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$6 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

.SUBCKT AOI211_X2 B A C2 C1 ZN NWELL|VDD VSS PWELL
M$1 \$12 B \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A \$12 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$11 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 \$5 B \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.055125P
+ PS=0.77U PD=0.805U
M$5 ZN C2 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.055125P AD=0.0441P
+ PS=0.805U PD=0.77U
M$6 \$5 C1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$7 ZN C1 \$5 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$8 \$5 C2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 ZN B VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$10 VSS A ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$11 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$12 VSS B ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0363125P
+ PS=0.555U PD=0.59U
M$13 \$13 C2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.0363125P AD=0.02905P
+ PS=0.59U PD=0.555U
M$14 ZN C1 \$13 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 \$14 C1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 VSS C2 \$14 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AOI211_X2

.SUBCKT MUX2_X1 A S B VSS NWELL|VDD Z PWELL
M$1 NWELL|VDD S \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.84U PD=0.455U
M$2 \$11 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P
+ AD=0.02205P PS=0.455U PD=0.455U
M$3 \$7 S \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P
+ PS=0.455U PD=0.455U
M$4 \$12 \$4 \$7 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P
+ PS=0.455U PD=0.455U
M$5 \$12 B NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.77U PD=0.455U
M$6 Z \$7 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P
+ PS=0.77U PD=1.47U
M$7 VSS S \$4 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$8 \$14 A VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$9 \$7 \$4 \$14 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$10 \$13 S \$7 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$11 VSS B \$13 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
M$12 Z \$7 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS MUX2_X1

.SUBCKT OR3_X1 A1 A2 A3 VSS NWELL|VDD ZN PWELL
M$1 \$11 A1 \$4 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P
+ PS=0.84U PD=0.455U
M$2 \$10 A2 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P
+ PS=0.455U PD=0.455U
M$3 \$10 A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.77U PD=0.455U
M$4 ZN \$4 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P
+ AD=0.06615P PS=0.77U PD=1.47U
M$5 VSS A1 \$4 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$6 \$4 A2 VSS PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U
+ PD=0.35U
M$7 VSS A3 \$4 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
M$8 ZN \$4 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OR3_X1

.SUBCKT AOI211_X1 C2 C1 B A VSS ZN NWELL|VDD PWELL
M$1 ZN C2 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$6 C1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$3 \$11 B \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 \$12 C2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$6 ZN C1 \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$7 VSS B ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$8 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI211_X1

.SUBCKT OAI211_X1 C2 C1 A B NWELL|VDD ZN VSS PWELL
M$1 \$11 C2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN C1 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 ZN B NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 ZN C2 \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$6 \$5 C1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$7 \$12 A \$5 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$8 VSS B \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OAI211_X1

.SUBCKT NAND3_X1 A3 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 ZN A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A2 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$4 \$10 A3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$5 \$9 A2 \$10 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$6 ZN A1 \$9 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NAND3_X1

.SUBCKT NOR3_X1 A3 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 \$10 A3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 \$9 A2 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 ZN A1 \$9 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$4 ZN A3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$5 VSS A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$6 ZN A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NOR3_X1

.SUBCKT OAI21_X1 B2 B1 A NWELL|VDD ZN VSS PWELL
M$1 \$10 B2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN B1 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 NWELL|VDD A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$4 ZN B2 \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$5 \$4 B1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$6 VSS A \$4 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS OAI21_X1

.SUBCKT NOR2_X4 A2 A1 ZN VSS NWELL|VDD PWELL
M$1 \$11 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN A1 \$11 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$10 A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 NWELL|VDD A2 \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$5 \$9 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$6 ZN A1 \$9 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$7 \$8 A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$8 NWELL|VDD A2 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$10 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 ZN A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 VSS A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$13 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$14 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 ZN A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$16 VSS A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NOR2_X4

.SUBCKT AND2_X1 A1 A2 NWELL|VDD VSS ZN PWELL
M$1 \$3 A1 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.84U PD=0.455U
M$2 \$3 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.77U PD=0.455U
M$3 ZN \$3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.033075P
+ AD=0.06615P PS=0.77U PD=1.47U
M$4 \$9 A1 \$3 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$5 VSS A2 \$9 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
M$6 ZN \$3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS AND2_X1

.SUBCKT NOR2_X1 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 \$8 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN A1 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$3 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$4 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NOR2_X1

.SUBCKT XNOR2_X1 A B NWELL|VDD VSS ZN PWELL
M$1 \$3 A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.033075P
+ AD=0.02205P PS=0.84U PD=0.455U
M$2 \$3 B NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.315U AS=0.0338625P
+ AD=0.02205P PS=0.775U PD=0.455U
M$3 ZN \$3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0338625P
+ AD=0.0441P PS=0.775U PD=0.77U
M$4 \$10 A ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$5 NWELL|VDD B \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$6 \$11 A \$3 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U
+ PD=0.35U
M$7 VSS B \$11 PWELL NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U
+ PD=0.56U
M$8 \$6 \$3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U
+ PD=0.555U
M$9 ZN A \$6 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$10 \$6 B ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS XNOR2_X1

.SUBCKT XOR2_X2 B A NWELL|VDD Z VSS PWELL
M$1 \$10 A \$3 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD B \$10 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$3 \$6 \$3 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P
+ PS=0.77U PD=0.77U
M$4 Z A \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$5 \$6 B Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$6 Z B \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$7 \$6 A Z NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$8 NWELL|VDD \$3 \$6 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$9 \$3 A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$10 VSS B \$3 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$11 Z \$3 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$12 \$12 A Z PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$13 VSS B \$12 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$14 \$11 B VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P
+ PS=0.555U PD=0.555U
M$15 Z A \$11 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$16 VSS \$3 Z PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS XOR2_X2

.SUBCKT NAND2_X1 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 ZN A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 NWELL|VDD A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$3 \$8 A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P
+ PS=1.04U PD=0.555U
M$4 ZN A1 \$8 PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NAND2_X1

.SUBCKT NOR2_X2 A2 A1 VSS NWELL|VDD ZN PWELL
M$1 \$9 A2 NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P
+ PS=1.47U PD=0.77U
M$2 ZN A1 \$9 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$3 \$8 A1 ZN NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U
+ PD=0.77U
M$4 NWELL|VDD A2 \$8 NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P
+ PS=0.77U PD=1.47U
M$5 ZN A2 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
M$6 VSS A1 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$7 ZN A1 VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
M$8 VSS A2 ZN PWELL NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P
+ PS=0.555U PD=1.04U
.ENDS NOR2_X2

.SUBCKT LOGIC0_X1 Z VSS NWELL|VDD PWELL
M$1 NWELL|VDD \$2 \$2 NWELL|VDD PMOS_VTL L=0.05U W=0.09U AS=0.00945P
+ AD=0.00945P PS=0.39U PD=0.39U
M$2 VSS \$2 Z PWELL NMOS_VTL L=0.05U W=0.09U AS=0.00945P AD=0.00945P PS=0.39U
+ PD=0.39U
.ENDS LOGIC0_X1

.SUBCKT INV_X1 A VSS NWELL|VDD ZN PWELL
M$1 ZN A NWELL|VDD NWELL|VDD PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P
+ PS=1.47U PD=1.47U
M$2 ZN A VSS PWELL NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

.SUBCKT TAPCELL_X1 VSS VDD PWELL NWELL
.ENDS TAPCELL_X1

.SUBCKT FILLCELL_X2 VSS NWELL|VDD PWELL
.ENDS FILLCELL_X2

.SUBCKT FILLCELL_X16 VSS NWELL|VDD PWELL
.ENDS FILLCELL_X16

.SUBCKT FILLCELL_X1 VSS NWELL|VDD PWELL
.ENDS FILLCELL_X1

.SUBCKT FILLCELL_X4 VSS NWELL|VDD PWELL
.ENDS FILLCELL_X4

.SUBCKT FILLCELL_X8 VSS NWELL|VDD PWELL
.ENDS FILLCELL_X8

.SUBCKT FILLCELL_X32 VSS NWELL|VDD PWELL
.ENDS FILLCELL_X32

.SUBCKT VIA_via1_7 \$1
.ENDS VIA_via1_7

.SUBCKT VIA_via3_2 \$1
.ENDS VIA_via3_2

.SUBCKT VIA_via5_0 \$1
.ENDS VIA_via5_0

.SUBCKT VIA_via4_0 \$1
.ENDS VIA_via4_0

.SUBCKT VIA_via5_6_940_1600_3_2_600_600 \$1
.ENDS VIA_via5_6_940_1600_3_2_600_600

.SUBCKT VIA_via6_7_940_1600_2_1_600_600 \$1
.ENDS VIA_via6_7_940_1600_2_1_600_600

.SUBCKT VIA_via1_2_940_340_1_3_300_300 \$1
.ENDS VIA_via1_2_940_340_1_3_300_300

.SUBCKT VIA_via2_3_940_340_1_3_320_320 \$1
.ENDS VIA_via2_3_940_340_1_3_320_320

.SUBCKT VIA_via3_4_940_340_1_3_320_320 \$1
.ENDS VIA_via3_4_940_340_1_3_320_320

.SUBCKT VIA_via7_8_940_1600_1_1_1680_1680 \$1
.ENDS VIA_via7_8_940_1600_1_1_1680_1680

.SUBCKT VIA_via8_9_940_1600_1_1_1680_1680 \$1
.ENDS VIA_via8_9_940_1600_1_1_1680_1680

.SUBCKT VIA_via9_10_1600_1600_1_1_3360_3360 \$1
.ENDS VIA_via9_10_1600_1600_1_1_3360_3360

.SUBCKT VIA_via4_5_940_1600_3_2_600_600 \$1
.ENDS VIA_via4_5_940_1600_3_2_600_600

.SUBCKT VIA_via4_5_940_960_2_2_600_600 \$1
.ENDS VIA_via4_5_940_960_2_2_600_600

.SUBCKT VIA_via5_6_940_960_2_2_600_600 \$1
.ENDS VIA_via5_6_940_960_2_2_600_600

.SUBCKT VIA_via6_7_940_960_1_1_600_600 \$1
.ENDS VIA_via6_7_940_960_1_1_600_600

.SUBCKT VIA_via7_8_1600_960_1_1_1680_1680 \$1
.ENDS VIA_via7_8_1600_960_1_1_1680_1680

.SUBCKT VIA_via2_5 \$1
.ENDS VIA_via2_5

.SUBCKT VIA_via1_4 \$1
.ENDS VIA_via1_4

.SUBCKT VIA_via8_9_1600_1600_1_1_1680_1680 \$1
.ENDS VIA_via8_9_1600_1600_1_1_1680_1680

.SUBCKT VIA_via9_10_1600_2400_1_1_3360_3360 \$1
.ENDS VIA_via9_10_1600_2400_1_1_3360_3360
