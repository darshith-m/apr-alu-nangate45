* Extracted by KLayout on : 19/02/2025 12:55

.SUBCKT spm
.ENDS spm
