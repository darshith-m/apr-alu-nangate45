module alu (clk,
    overflow_flag,
    rst_n,
    zero_flag,
    a,
    b,
    opcode,
    result);
 input clk;
 output overflow_flag;
 input rst_n;
 output zero_flag;
 input [7:0] a;
 input [7:0] b;
 input [3:0] opcode;
 output [7:0] result;

 wire clknet_0_clk;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;

 INV_X1 _239_ (.A(a[1]),
    .ZN(_162_));
 INV_X2 _240_ (.A(net44),
    .ZN(_163_));
 INV_X1 _241_ (.A(net107),
    .ZN(_164_));
 INV_X2 _242_ (.A(net45),
    .ZN(_165_));
 INV_X1 _243_ (.A(a[5]),
    .ZN(_166_));
 INV_X1 _244_ (.A(a[6]),
    .ZN(_167_));
 INV_X2 _245_ (.A(b[2]),
    .ZN(_168_));
 INV_X1 _246_ (.A(net74),
    .ZN(_169_));
 INV_X1 _247_ (.A(b[4]),
    .ZN(_170_));
 INV_X1 _248_ (.A(b[5]),
    .ZN(_171_));
 INV_X1 _249_ (.A(net65),
    .ZN(_172_));
 INV_X1 _250_ (.A(net80),
    .ZN(_173_));
 INV_X1 _251_ (.A(opcode[3]),
    .ZN(_174_));
 INV_X1 _252_ (.A(net50),
    .ZN(_175_));
 NOR2_X2 _253_ (.A1(net51),
    .A2(net49),
    .ZN(_176_));
 INV_X1 _254_ (.A(_176_),
    .ZN(_177_));
 NAND2_X1 _255_ (.A1(net48),
    .A2(_172_),
    .ZN(_178_));
 NAND2_X1 _256_ (.A1(net48),
    .A2(net65),
    .ZN(_179_));
 XOR2_X2 _257_ (.A(net48),
    .B(net65),
    .Z(_180_));
 XNOR2_X1 _258_ (.A(net48),
    .B(net65),
    .ZN(_181_));
 NOR2_X1 _259_ (.A1(_167_),
    .A2(net104),
    .ZN(_182_));
 OR2_X1 _260_ (.A1(a[6]),
    .A2(b[6]),
    .ZN(_183_));
 NAND2_X2 _261_ (.A1(a[6]),
    .A2(net104),
    .ZN(_184_));
 AND2_X1 _262_ (.A1(_183_),
    .A2(_184_),
    .ZN(_185_));
 NAND2_X1 _263_ (.A1(_183_),
    .A2(_184_),
    .ZN(_186_));
 NOR2_X2 _264_ (.A1(_164_),
    .A2(b[3]),
    .ZN(_187_));
 AND2_X1 _265_ (.A1(net107),
    .A2(b[3]),
    .ZN(_188_));
 NOR2_X2 _266_ (.A1(net107),
    .A2(b[3]),
    .ZN(_189_));
 INV_X1 _267_ (.A(net108),
    .ZN(_190_));
 NOR2_X4 _268_ (.A1(net41),
    .A2(net108),
    .ZN(_191_));
 NAND2_X1 _269_ (.A1(a[2]),
    .A2(_168_),
    .ZN(_192_));
 OR2_X1 _270_ (.A1(net138),
    .A2(b[2]),
    .ZN(_193_));
 NAND2_X1 _271_ (.A1(a[2]),
    .A2(b[2]),
    .ZN(_194_));
 AND2_X1 _272_ (.A1(_193_),
    .A2(_194_),
    .ZN(_195_));
 NAND2_X2 _273_ (.A1(_193_),
    .A2(_194_),
    .ZN(_196_));
 AND2_X1 _274_ (.A1(a[1]),
    .A2(net45),
    .ZN(_197_));
 XOR2_X2 _275_ (.A(a[1]),
    .B(net45),
    .Z(_198_));
 AOI21_X2 _276_ (.A(_198_),
    .B1(_169_),
    .B2(net43),
    .ZN(_199_));
 NOR2_X1 _277_ (.A1(_162_),
    .A2(net45),
    .ZN(_200_));
 OAI21_X2 _278_ (.A(_196_),
    .B1(_199_),
    .B2(_200_),
    .ZN(_201_));
 AOI21_X4 _279_ (.A(_191_),
    .B1(_192_),
    .B2(_201_),
    .ZN(_202_));
 NOR2_X1 _280_ (.A1(_187_),
    .A2(_202_),
    .ZN(_203_));
 NOR2_X1 _281_ (.A1(_166_),
    .A2(_171_),
    .ZN(_204_));
 XOR2_X2 _282_ (.A(a[5]),
    .B(b[5]),
    .Z(_205_));
 XNOR2_X2 _283_ (.A(a[5]),
    .B(b[5]),
    .ZN(_206_));
 NAND2_X1 _284_ (.A1(net47),
    .A2(net114),
    .ZN(_207_));
 XOR2_X2 _285_ (.A(net47),
    .B(net114),
    .Z(_208_));
 XNOR2_X2 _286_ (.A(net47),
    .B(net114),
    .ZN(_209_));
 NAND2_X1 _287_ (.A1(_206_),
    .A2(_209_),
    .ZN(_210_));
 OAI211_X2 _288_ (.A(_206_),
    .B(_209_),
    .C1(_187_),
    .C2(_202_),
    .ZN(_211_));
 NAND2_X1 _289_ (.A1(net91),
    .A2(_170_),
    .ZN(_212_));
 NOR2_X1 _290_ (.A1(_205_),
    .A2(net92),
    .ZN(_213_));
 AOI21_X2 _291_ (.A(_213_),
    .B1(_171_),
    .B2(net141),
    .ZN(_214_));
 AOI21_X2 _292_ (.A(net40),
    .B1(_211_),
    .B2(_214_),
    .ZN(_215_));
 NOR2_X1 _293_ (.A1(net105),
    .A2(_215_),
    .ZN(_216_));
 OAI21_X1 _294_ (.A(_181_),
    .B1(_182_),
    .B2(_215_),
    .ZN(_217_));
 AND2_X1 _295_ (.A1(_178_),
    .A2(_217_),
    .ZN(_218_));
 NAND2_X1 _296_ (.A1(_178_),
    .A2(_217_),
    .ZN(_219_));
 NAND2_X4 _297_ (.A1(_174_),
    .A2(net69),
    .ZN(_220_));
 NAND2_X2 _298_ (.A1(net80),
    .A2(opcode[1]),
    .ZN(_221_));
 NOR2_X1 _299_ (.A1(net70),
    .A2(_221_),
    .ZN(_222_));
 NOR2_X1 _300_ (.A1(net43),
    .A2(_169_),
    .ZN(_223_));
 AND2_X1 _301_ (.A1(net43),
    .A2(net74),
    .ZN(_224_));
 NAND2_X1 _302_ (.A1(net43),
    .A2(net74),
    .ZN(_225_));
 NAND2_X1 _303_ (.A1(_163_),
    .A2(_169_),
    .ZN(_226_));
 NOR2_X1 _304_ (.A1(_191_),
    .A2(_223_),
    .ZN(_227_));
 NOR3_X1 _305_ (.A1(_180_),
    .A2(net40),
    .A3(_195_),
    .ZN(_228_));
 NAND3_X1 _306_ (.A1(_199_),
    .A2(_227_),
    .A3(_228_),
    .ZN(_011_));
 OAI21_X1 _307_ (.A(net71),
    .B1(_011_),
    .B2(_210_),
    .ZN(_012_));
 INV_X1 _308_ (.A(_012_),
    .ZN(_013_));
 OR2_X4 _309_ (.A1(net144),
    .A2(net69),
    .ZN(_014_));
 NOR2_X2 _310_ (.A1(opcode[1]),
    .A2(_014_),
    .ZN(_015_));
 NOR2_X2 _311_ (.A1(opcode[1]),
    .A2(_220_),
    .ZN(_016_));
 NOR3_X4 _312_ (.A1(net80),
    .A2(opcode[1]),
    .A3(net70),
    .ZN(_017_));
 OAI211_X1 _313_ (.A(net75),
    .B(_226_),
    .C1(_015_),
    .C2(_017_),
    .ZN(_018_));
 NOR2_X4 _314_ (.A1(_221_),
    .A2(_014_),
    .ZN(_019_));
 NAND2_X1 _315_ (.A1(_226_),
    .A2(_019_),
    .ZN(_020_));
 NAND2_X2 _316_ (.A1(_173_),
    .A2(opcode[1]),
    .ZN(_021_));
 OR2_X2 _317_ (.A1(_014_),
    .A2(_021_),
    .ZN(_022_));
 INV_X1 _318_ (.A(_022_),
    .ZN(_023_));
 OAI211_X1 _319_ (.A(net76),
    .B(_020_),
    .C1(_022_),
    .C2(net75),
    .ZN(_024_));
 AOI211_X1 _320_ (.A(net45),
    .B(_223_),
    .C1(a[1]),
    .C2(net43),
    .ZN(_025_));
 AND2_X1 _321_ (.A1(a[2]),
    .A2(_163_),
    .ZN(_026_));
 NOR2_X1 _322_ (.A1(_163_),
    .A2(_164_),
    .ZN(_027_));
 NOR2_X1 _323_ (.A1(_026_),
    .A2(_027_),
    .ZN(_028_));
 NOR3_X4 _324_ (.A1(b[2]),
    .A2(net70),
    .A3(_021_),
    .ZN(_029_));
 OR3_X2 _325_ (.A1(b[2]),
    .A2(_220_),
    .A3(_021_),
    .ZN(_030_));
 AOI211_X1 _326_ (.A(_025_),
    .B(_030_),
    .C1(_028_),
    .C2(net45),
    .ZN(_031_));
 NOR3_X1 _327_ (.A1(_168_),
    .A2(net70),
    .A3(_021_),
    .ZN(_032_));
 OR3_X1 _328_ (.A1(_168_),
    .A2(_220_),
    .A3(_021_),
    .ZN(_033_));
 MUX2_X1 _329_ (.A(net47),
    .B(a[5]),
    .S(net44),
    .Z(_034_));
 NOR2_X1 _330_ (.A1(net44),
    .A2(_167_),
    .ZN(_035_));
 AOI21_X2 _331_ (.A(_035_),
    .B1(net48),
    .B2(net44),
    .ZN(_036_));
 NOR2_X1 _332_ (.A1(net42),
    .A2(_034_),
    .ZN(_037_));
 AOI211_X1 _333_ (.A(_033_),
    .B(_037_),
    .C1(_036_),
    .C2(net32),
    .ZN(_038_));
 NOR3_X1 _334_ (.A1(net43),
    .A2(net45),
    .A3(_169_),
    .ZN(_039_));
 NAND2_X1 _335_ (.A1(net80),
    .A2(_016_),
    .ZN(_040_));
 NOR2_X2 _336_ (.A1(b[2]),
    .A2(_040_),
    .ZN(_041_));
 NAND3_X4 _337_ (.A1(_168_),
    .A2(net80),
    .A3(_016_),
    .ZN(_042_));
 AND2_X1 _338_ (.A1(_039_),
    .A2(_041_),
    .ZN(_043_));
 OR3_X1 _339_ (.A1(_031_),
    .A2(_038_),
    .A3(_043_),
    .ZN(_044_));
 AOI211_X2 _340_ (.A(net77),
    .B(_044_),
    .C1(_219_),
    .C2(_013_),
    .ZN(_045_));
 AOI21_X1 _341_ (.A(_176_),
    .B1(net78),
    .B2(net27),
    .ZN(_001_));
 AOI211_X1 _342_ (.A(_221_),
    .B(_014_),
    .C1(_162_),
    .C2(_165_),
    .ZN(_046_));
 AOI221_X1 _343_ (.A(_046_),
    .B1(_017_),
    .B2(_198_),
    .C1(_197_),
    .C2(_023_),
    .ZN(_047_));
 NOR2_X1 _344_ (.A1(net44),
    .A2(_166_),
    .ZN(_048_));
 AOI21_X2 _345_ (.A(_048_),
    .B1(a[6]),
    .B2(net35),
    .ZN(_049_));
 NAND2_X1 _346_ (.A1(_163_),
    .A2(net48),
    .ZN(_050_));
 NAND3_X1 _347_ (.A1(_163_),
    .A2(net42),
    .A3(net48),
    .ZN(_051_));
 OAI21_X2 _348_ (.A(_051_),
    .B1(_049_),
    .B2(net42),
    .ZN(_052_));
 NAND2_X2 _349_ (.A1(net80),
    .A2(_015_),
    .ZN(_053_));
 NAND3_X1 _350_ (.A1(net43),
    .A2(_169_),
    .A3(_198_),
    .ZN(_054_));
 NOR2_X1 _351_ (.A1(_199_),
    .A2(_053_),
    .ZN(_055_));
 NOR3_X1 _352_ (.A1(net137),
    .A2(opcode[1]),
    .A3(_014_),
    .ZN(_056_));
 NAND2_X2 _353_ (.A1(_173_),
    .A2(_015_),
    .ZN(_057_));
 XNOR2_X1 _354_ (.A(_198_),
    .B(_225_),
    .ZN(_058_));
 NOR2_X1 _355_ (.A1(_162_),
    .A2(net43),
    .ZN(_059_));
 NOR2_X1 _356_ (.A1(_224_),
    .A2(_059_),
    .ZN(_060_));
 NOR3_X1 _357_ (.A1(net32),
    .A2(_042_),
    .A3(_060_),
    .ZN(_061_));
 AOI21_X1 _358_ (.A(_059_),
    .B1(net37),
    .B2(a[2]),
    .ZN(_062_));
 MUX2_X1 _359_ (.A(net107),
    .B(net47),
    .S(net44),
    .Z(_063_));
 OAI21_X1 _360_ (.A(_029_),
    .B1(_063_),
    .B2(_165_),
    .ZN(_064_));
 AOI21_X1 _361_ (.A(_064_),
    .B1(_062_),
    .B2(_165_),
    .ZN(_065_));
 AOI21_X1 _362_ (.A(_061_),
    .B1(_052_),
    .B2(_032_),
    .ZN(_066_));
 AOI221_X1 _363_ (.A(_065_),
    .B1(_058_),
    .B2(_056_),
    .C1(_054_),
    .C2(_055_),
    .ZN(_067_));
 NAND3_X1 _364_ (.A1(_047_),
    .A2(_066_),
    .A3(_067_),
    .ZN(_068_));
 AOI21_X1 _365_ (.A(_068_),
    .B1(net71),
    .B2(_218_),
    .ZN(_069_));
 AOI21_X1 _366_ (.A(_176_),
    .B1(net72),
    .B2(net27),
    .ZN(_002_));
 OR3_X1 _367_ (.A1(_196_),
    .A2(_199_),
    .A3(_200_),
    .ZN(_070_));
 NAND4_X1 _368_ (.A1(net80),
    .A2(_201_),
    .A3(_015_),
    .A4(_070_),
    .ZN(_071_));
 AOI21_X2 _369_ (.A(_197_),
    .B1(_198_),
    .B2(_224_),
    .ZN(_072_));
 OAI211_X1 _370_ (.A(_173_),
    .B(_015_),
    .C1(_072_),
    .C2(_196_),
    .ZN(_073_));
 AOI21_X1 _371_ (.A(_073_),
    .B1(_072_),
    .B2(_196_),
    .ZN(_074_));
 OR3_X1 _372_ (.A1(net32),
    .A2(_033_),
    .A3(_036_),
    .ZN(_075_));
 AOI21_X2 _373_ (.A(_026_),
    .B1(net44),
    .B2(a[1]),
    .ZN(_076_));
 NAND2_X1 _374_ (.A1(net45),
    .A2(_223_),
    .ZN(_077_));
 OAI21_X2 _375_ (.A(_077_),
    .B1(_076_),
    .B2(net46),
    .ZN(_078_));
 NAND2_X1 _376_ (.A1(net46),
    .A2(_034_),
    .ZN(_079_));
 OAI21_X1 _377_ (.A(_079_),
    .B1(_028_),
    .B2(net42),
    .ZN(_080_));
 AOI221_X1 _378_ (.A(_074_),
    .B1(_078_),
    .B2(_041_),
    .C1(_019_),
    .C2(_193_),
    .ZN(_081_));
 OAI211_X1 _379_ (.A(net49),
    .B(_075_),
    .C1(_022_),
    .C2(_194_),
    .ZN(_082_));
 AOI221_X2 _380_ (.A(_082_),
    .B1(_080_),
    .B2(_029_),
    .C1(_195_),
    .C2(_017_),
    .ZN(_083_));
 NAND3_X1 _381_ (.A1(net81),
    .A2(net139),
    .A3(_083_),
    .ZN(_084_));
 AND2_X1 _382_ (.A1(_177_),
    .A2(net82),
    .ZN(_003_));
 OAI21_X1 _383_ (.A(_194_),
    .B1(_196_),
    .B2(_072_),
    .ZN(_085_));
 XNOR2_X1 _384_ (.A(_191_),
    .B(_085_),
    .ZN(_086_));
 NOR2_X1 _385_ (.A1(_057_),
    .A2(_086_),
    .ZN(_087_));
 AND3_X1 _386_ (.A1(_191_),
    .A2(_192_),
    .A3(_201_),
    .ZN(_088_));
 NOR3_X1 _387_ (.A1(_202_),
    .A2(_053_),
    .A3(_088_),
    .ZN(_089_));
 NOR3_X1 _388_ (.A1(net46),
    .A2(_033_),
    .A3(_050_),
    .ZN(_090_));
 MUX2_X1 _389_ (.A(a[3]),
    .B(a[2]),
    .S(net44),
    .Z(_091_));
 NAND2_X1 _390_ (.A1(_165_),
    .A2(_091_),
    .ZN(_092_));
 OAI21_X1 _391_ (.A(_092_),
    .B1(_060_),
    .B2(_165_),
    .ZN(_093_));
 AOI21_X1 _392_ (.A(_030_),
    .B1(_049_),
    .B2(net42),
    .ZN(_094_));
 OAI21_X1 _393_ (.A(_094_),
    .B1(_063_),
    .B2(net42),
    .ZN(_095_));
 AOI221_X1 _394_ (.A(_090_),
    .B1(_093_),
    .B2(_041_),
    .C1(_023_),
    .C2(net41),
    .ZN(_096_));
 AOI22_X1 _395_ (.A1(_191_),
    .A2(_017_),
    .B1(_019_),
    .B2(net109),
    .ZN(_097_));
 NAND3_X1 _396_ (.A1(_095_),
    .A2(_096_),
    .A3(net110),
    .ZN(_098_));
 OR3_X1 _397_ (.A1(_087_),
    .A2(_089_),
    .A3(net111),
    .ZN(_099_));
 MUX2_X1 _398_ (.A(net52),
    .B(net112),
    .S(net27),
    .Z(_004_));
 NOR2_X1 _399_ (.A1(_203_),
    .A2(_208_),
    .ZN(_100_));
 NOR3_X1 _400_ (.A1(_187_),
    .A2(_202_),
    .A3(_209_),
    .ZN(_101_));
 OR3_X1 _401_ (.A1(_053_),
    .A2(_100_),
    .A3(_101_),
    .ZN(_102_));
 AOI21_X1 _402_ (.A(net41),
    .B1(_191_),
    .B2(_085_),
    .ZN(_103_));
 XNOR2_X1 _403_ (.A(_209_),
    .B(_103_),
    .ZN(_104_));
 AOI21_X1 _404_ (.A(_027_),
    .B1(net47),
    .B2(_163_),
    .ZN(_105_));
 AND2_X1 _405_ (.A1(_165_),
    .A2(_105_),
    .ZN(_106_));
 AOI211_X2 _406_ (.A(_042_),
    .B(_106_),
    .C1(_076_),
    .C2(net46),
    .ZN(_107_));
 OAI21_X1 _407_ (.A(_019_),
    .B1(net114),
    .B2(net47),
    .ZN(_108_));
 OAI21_X1 _408_ (.A(_108_),
    .B1(_022_),
    .B2(_207_),
    .ZN(_109_));
 AOI211_X1 _409_ (.A(_107_),
    .B(_109_),
    .C1(_208_),
    .C2(_017_),
    .ZN(_110_));
 AOI211_X1 _410_ (.A(_030_),
    .B(_037_),
    .C1(_036_),
    .C2(net46),
    .ZN(_111_));
 NOR2_X1 _411_ (.A1(_168_),
    .A2(_040_),
    .ZN(_112_));
 AOI21_X1 _412_ (.A(_111_),
    .B1(_112_),
    .B2(_039_),
    .ZN(_113_));
 AND2_X1 _413_ (.A1(net115),
    .A2(_113_),
    .ZN(_114_));
 OAI211_X1 _414_ (.A(_102_),
    .B(_114_),
    .C1(_104_),
    .C2(_057_),
    .ZN(_115_));
 MUX2_X1 _415_ (.A(net53),
    .B(net116),
    .S(net27),
    .Z(_005_));
 OAI21_X1 _416_ (.A(_207_),
    .B1(_209_),
    .B2(_103_),
    .ZN(_116_));
 XNOR2_X1 _417_ (.A(_205_),
    .B(_116_),
    .ZN(_117_));
 NAND2_X1 _418_ (.A1(_205_),
    .A2(net92),
    .ZN(_118_));
 NOR2_X1 _419_ (.A1(_213_),
    .A2(_053_),
    .ZN(_119_));
 OAI211_X1 _420_ (.A(_211_),
    .B(_119_),
    .C1(net93),
    .C2(_100_),
    .ZN(_120_));
 AOI211_X2 _421_ (.A(_221_),
    .B(_014_),
    .C1(_166_),
    .C2(_171_),
    .ZN(_121_));
 AOI221_X2 _422_ (.A(_121_),
    .B1(_017_),
    .B2(_205_),
    .C1(_204_),
    .C2(_023_),
    .ZN(_122_));
 OR4_X1 _423_ (.A1(net32),
    .A2(_168_),
    .A3(_040_),
    .A4(_060_),
    .ZN(_123_));
 NAND2_X1 _424_ (.A1(_122_),
    .A2(_123_),
    .ZN(_124_));
 AOI21_X2 _425_ (.A(_048_),
    .B1(net47),
    .B2(net35),
    .ZN(_125_));
 NOR2_X1 _426_ (.A1(_165_),
    .A2(_091_),
    .ZN(_126_));
 AOI211_X2 _427_ (.A(_042_),
    .B(_126_),
    .C1(_125_),
    .C2(_165_),
    .ZN(_127_));
 AOI211_X2 _428_ (.A(_124_),
    .B(_127_),
    .C1(_029_),
    .C2(_052_),
    .ZN(_128_));
 OAI211_X1 _429_ (.A(net94),
    .B(_128_),
    .C1(_057_),
    .C2(_117_),
    .ZN(_129_));
 INV_X1 _430_ (.A(net95),
    .ZN(_130_));
 AOI21_X1 _431_ (.A(_176_),
    .B1(net96),
    .B2(net27),
    .ZN(_006_));
 AOI21_X1 _432_ (.A(_204_),
    .B1(_205_),
    .B2(_116_),
    .ZN(_131_));
 OR2_X1 _433_ (.A1(_186_),
    .A2(_131_),
    .ZN(_132_));
 AOI21_X1 _434_ (.A(_057_),
    .B1(_131_),
    .B2(_186_),
    .ZN(_133_));
 NAND3_X1 _435_ (.A1(net40),
    .A2(_211_),
    .A3(net142),
    .ZN(_134_));
 NOR2_X1 _436_ (.A1(_215_),
    .A2(_053_),
    .ZN(_135_));
 NOR3_X1 _437_ (.A1(net46),
    .A2(_030_),
    .A3(_036_),
    .ZN(_136_));
 NOR2_X1 _438_ (.A1(_184_),
    .A2(_022_),
    .ZN(_137_));
 AOI21_X1 _439_ (.A(_136_),
    .B1(_017_),
    .B2(net40),
    .ZN(_138_));
 MUX2_X1 _440_ (.A(a[6]),
    .B(a[5]),
    .S(net35),
    .Z(_139_));
 NAND2_X1 _441_ (.A1(net42),
    .A2(_105_),
    .ZN(_140_));
 OAI211_X1 _442_ (.A(_041_),
    .B(_140_),
    .C1(_139_),
    .C2(net99),
    .ZN(_141_));
 AOI221_X2 _443_ (.A(_137_),
    .B1(_112_),
    .B2(_078_),
    .C1(_183_),
    .C2(_019_),
    .ZN(_142_));
 NAND3_X1 _444_ (.A1(_138_),
    .A2(net100),
    .A3(_142_),
    .ZN(_143_));
 AOI221_X2 _445_ (.A(net101),
    .B1(_135_),
    .B2(_134_),
    .C1(_132_),
    .C2(_133_),
    .ZN(_144_));
 AOI21_X1 _446_ (.A(_176_),
    .B1(net102),
    .B2(net27),
    .ZN(_007_));
 AOI21_X1 _447_ (.A(_181_),
    .B1(_184_),
    .B2(_132_),
    .ZN(_145_));
 AND3_X1 _448_ (.A1(_181_),
    .A2(_184_),
    .A3(_132_),
    .ZN(_146_));
 OR2_X1 _449_ (.A1(_057_),
    .A2(_145_),
    .ZN(_147_));
 XNOR2_X1 _450_ (.A(_180_),
    .B(_216_),
    .ZN(_148_));
 AOI211_X1 _451_ (.A(net46),
    .B(_050_),
    .C1(_042_),
    .C2(_030_),
    .ZN(_149_));
 AOI21_X1 _452_ (.A(net42),
    .B1(a[6]),
    .B2(net35),
    .ZN(_150_));
 AOI211_X1 _453_ (.A(_042_),
    .B(_150_),
    .C1(_125_),
    .C2(net33),
    .ZN(_151_));
 AND2_X1 _454_ (.A1(_093_),
    .A2(_112_),
    .ZN(_152_));
 OAI21_X1 _455_ (.A(_019_),
    .B1(net65),
    .B2(net84),
    .ZN(_153_));
 OAI21_X1 _456_ (.A(net85),
    .B1(_022_),
    .B2(_179_),
    .ZN(_154_));
 OR3_X1 _457_ (.A1(_149_),
    .A2(_151_),
    .A3(net86),
    .ZN(_155_));
 AOI211_X2 _458_ (.A(_152_),
    .B(net87),
    .C1(_180_),
    .C2(_017_),
    .ZN(_156_));
 OAI221_X1 _459_ (.A(net88),
    .B1(_147_),
    .B2(_146_),
    .C1(_053_),
    .C2(_148_),
    .ZN(_157_));
 MUX2_X1 _460_ (.A(net54),
    .B(net89),
    .S(net27),
    .Z(_008_));
 NOR4_X1 _461_ (.A1(net82),
    .A2(net112),
    .A3(_115_),
    .A4(net95),
    .ZN(_158_));
 NAND4_X1 _462_ (.A1(net78),
    .A2(net72),
    .A3(net102),
    .A4(_158_),
    .ZN(_159_));
 OAI22_X1 _463_ (.A1(_175_),
    .A2(net27),
    .B1(net89),
    .B2(_159_),
    .ZN(_009_));
 AOI21_X1 _464_ (.A(_145_),
    .B1(net65),
    .B2(net48),
    .ZN(_160_));
 OAI221_X1 _465_ (.A(net49),
    .B1(_219_),
    .B2(_053_),
    .C1(_057_),
    .C2(net66),
    .ZN(_161_));
 AND2_X1 _466_ (.A1(_177_),
    .A2(net67),
    .ZN(_010_));
 DFF_X2 _467_ (.D(net79),
    .CK(clknet_1_1__leaf_clk),
    .Q(net61),
    .QN(_238_));
 DFF_X2 _468_ (.D(net73),
    .CK(clknet_1_1__leaf_clk),
    .Q(net62),
    .QN(_237_));
 DFF_X2 _469_ (.D(net83),
    .CK(clknet_1_1__leaf_clk),
    .Q(net63),
    .QN(_236_));
 DFF_X2 _470_ (.D(net113),
    .CK(clknet_1_0__leaf_clk),
    .Q(net57),
    .QN(_235_));
 DFF_X2 _471_ (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net55),
    .QN(_234_));
 DFF_X2 _472_ (.D(net97),
    .CK(clknet_1_0__leaf_clk),
    .Q(net58),
    .QN(_233_));
 DFF_X2 _473_ (.D(net103),
    .CK(clknet_1_0__leaf_clk),
    .Q(net60),
    .QN(_232_));
 DFF_X2 _474_ (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net59),
    .QN(_231_));
 DFF_X2 _475_ (.D(net90),
    .CK(clknet_1_0__leaf_clk),
    .Q(net56),
    .QN(_230_));
 DFF_X2 _476_ (.D(net68),
    .CK(clknet_1_1__leaf_clk),
    .Q(net64),
    .QN(_229_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 TAPCELL_X1 TAP_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 TAP_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 TAP_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 TAP_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 TAP_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 TAP_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 TAP_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 TAP_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 TAP_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 TAP_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 TAP_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 TAP_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 TAP_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 TAP_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 TAP_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 TAP_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 TAP_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 TAP_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 TAP_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 TAP_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 TAP_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 TAP_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 TAP_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 TAP_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 TAP_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 TAP_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 TAP_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 TAP_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 TAP_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 TAP_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 TAP_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 TAP_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 TAP_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 TAP_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 TAP_EDGE_ROW_0_Left_34 ();
 TAPCELL_X1 TAP_EDGE_ROW_1_Left_35 ();
 TAPCELL_X1 TAP_EDGE_ROW_2_Left_36 ();
 TAPCELL_X1 TAP_EDGE_ROW_3_Left_37 ();
 TAPCELL_X1 TAP_EDGE_ROW_4_Left_38 ();
 TAPCELL_X1 TAP_EDGE_ROW_5_Left_39 ();
 TAPCELL_X1 TAP_EDGE_ROW_6_Left_40 ();
 TAPCELL_X1 TAP_EDGE_ROW_7_Left_41 ();
 TAPCELL_X1 TAP_EDGE_ROW_8_Left_42 ();
 TAPCELL_X1 TAP_EDGE_ROW_9_Left_43 ();
 TAPCELL_X1 TAP_EDGE_ROW_10_Left_44 ();
 TAPCELL_X1 TAP_EDGE_ROW_11_Left_45 ();
 TAPCELL_X1 TAP_EDGE_ROW_12_Left_46 ();
 TAPCELL_X1 TAP_EDGE_ROW_13_Left_47 ();
 TAPCELL_X1 TAP_EDGE_ROW_14_Left_48 ();
 TAPCELL_X1 TAP_EDGE_ROW_15_Left_49 ();
 TAPCELL_X1 TAP_EDGE_ROW_16_Left_50 ();
 TAPCELL_X1 TAP_EDGE_ROW_17_Left_51 ();
 TAPCELL_X1 TAP_EDGE_ROW_18_Left_52 ();
 TAPCELL_X1 TAP_EDGE_ROW_19_Left_53 ();
 TAPCELL_X1 TAP_EDGE_ROW_20_Left_54 ();
 TAPCELL_X1 TAP_EDGE_ROW_21_Left_55 ();
 TAPCELL_X1 TAP_EDGE_ROW_22_Left_56 ();
 TAPCELL_X1 TAP_EDGE_ROW_23_Left_57 ();
 TAPCELL_X1 TAP_EDGE_ROW_24_Left_58 ();
 TAPCELL_X1 TAP_EDGE_ROW_25_Left_59 ();
 TAPCELL_X1 TAP_EDGE_ROW_26_Left_60 ();
 TAPCELL_X1 TAP_EDGE_ROW_27_Left_61 ();
 TAPCELL_X1 TAP_EDGE_ROW_28_Left_62 ();
 TAPCELL_X1 TAP_EDGE_ROW_29_Left_63 ();
 TAPCELL_X1 TAP_EDGE_ROW_30_Left_64 ();
 TAPCELL_X1 TAP_EDGE_ROW_31_Left_65 ();
 TAPCELL_X1 TAP_EDGE_ROW_32_Left_66 ();
 TAPCELL_X1 TAP_EDGE_ROW_33_Left_67 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_68 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_69 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_70 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_71 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_72 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_73 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_74 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_75 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_76 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_77 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_78 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_79 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_80 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_81 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_82 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_83 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_84 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_85 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_86 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_87 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_88 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_89 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_90 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_91 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_92 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_93 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_94 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_95 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_96 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_97 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_98 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_99 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_121 ();
 BUF_X2 fanout27 (.A(net49),
    .Z(net27));
 BUF_X1 fanout28 (.A(rst_n),
    .Z(net28));
 BUF_X2 fanout29 (.A(net46),
    .Z(net29));
 BUF_X1 fanout30 (.A(net33),
    .Z(net30));
 BUF_X1 fanout31 (.A(net33),
    .Z(net31));
 BUF_X1 fanout32 (.A(net33),
    .Z(net32));
 BUF_X1 fanout33 (.A(net98),
    .Z(net33));
 BUF_X1 fanout34 (.A(net37),
    .Z(net34));
 CLKBUF_X2 fanout35 (.A(net37),
    .Z(net35));
 BUF_X2 fanout36 (.A(net37),
    .Z(net36));
 BUF_X1 fanout37 (.A(b[0]),
    .Z(net37));
 BUF_X1 fanout38 (.A(net84),
    .Z(net38));
 BUF_X1 fanout39 (.A(net91),
    .Z(net39));
 BUF_X2 gain40 (.A(_185_),
    .Z(net40));
 BUF_X2 gain41 (.A(_188_),
    .Z(net41));
 BUF_X4 gain42 (.A(net29),
    .Z(net42));
 BUF_X4 gain43 (.A(net36),
    .Z(net43));
 BUF_X4 gain44 (.A(net34),
    .Z(net44));
 BUF_X4 gain45 (.A(net31),
    .Z(net45));
 BUF_X4 gain46 (.A(net30),
    .Z(net46));
 BUF_X4 gain47 (.A(net39),
    .Z(net47));
 BUF_X4 gain48 (.A(net38),
    .Z(net48));
 BUF_X2 gain49 (.A(net28),
    .Z(net49));
 LOGIC0_X1 _252__50 (.Z(net50));
 LOGIC0_X1 _253__51 (.Z(net51));
 LOGIC0_X1 _398__52 (.Z(net52));
 LOGIC0_X1 _415__53 (.Z(net53));
 LOGIC0_X1 _460__54 (.Z(net54));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 CLKBUF_X1 hold55 (.A(net117),
    .Z(net118));
 CLKBUF_X1 hold56 (.A(net119),
    .Z(net120));
 CLKBUF_X1 hold57 (.A(net121),
    .Z(net122));
 CLKBUF_X1 hold58 (.A(net123),
    .Z(net124));
 CLKBUF_X1 hold59 (.A(net125),
    .Z(net126));
 CLKBUF_X1 hold60 (.A(net127),
    .Z(net128));
 CLKBUF_X1 hold61 (.A(net129),
    .Z(net130));
 CLKBUF_X1 hold62 (.A(net131),
    .Z(net132));
 CLKBUF_X1 hold63 (.A(net133),
    .Z(net134));
 CLKBUF_X1 hold64 (.A(net135),
    .Z(net136));
 CLKBUF_X1 hold65 (.A(b[7]),
    .Z(net65));
 CLKBUF_X1 hold66 (.A(_160_),
    .Z(net66));
 CLKBUF_X1 hold67 (.A(_161_),
    .Z(net67));
 CLKBUF_X1 hold68 (.A(_010_),
    .Z(net68));
 CLKBUF_X1 hold69 (.A(opcode[2]),
    .Z(net69));
 CLKBUF_X1 hold70 (.A(_220_),
    .Z(net70));
 CLKBUF_X1 hold71 (.A(_222_),
    .Z(net71));
 CLKBUF_X1 hold72 (.A(_069_),
    .Z(net72));
 CLKBUF_X1 hold73 (.A(_002_),
    .Z(net73));
 CLKBUF_X1 hold74 (.A(a[0]),
    .Z(net74));
 CLKBUF_X1 hold75 (.A(_225_),
    .Z(net75));
 CLKBUF_X1 hold76 (.A(_018_),
    .Z(net76));
 CLKBUF_X1 hold77 (.A(_024_),
    .Z(net77));
 CLKBUF_X1 hold78 (.A(_045_),
    .Z(net78));
 CLKBUF_X1 hold79 (.A(_001_),
    .Z(net79));
 CLKBUF_X1 hold80 (.A(opcode[0]),
    .Z(net80));
 CLKBUF_X1 hold81 (.A(_071_),
    .Z(net81));
 CLKBUF_X1 hold82 (.A(net140),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(_003_),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(a[7]),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(_153_),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(_154_),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(_155_),
    .Z(net87));
 CLKBUF_X1 hold88 (.A(_156_),
    .Z(net88));
 CLKBUF_X1 hold89 (.A(net106),
    .Z(net89));
 CLKBUF_X1 hold90 (.A(_009_),
    .Z(net90));
 CLKBUF_X1 hold91 (.A(a[4]),
    .Z(net91));
 CLKBUF_X1 hold92 (.A(_212_),
    .Z(net92));
 CLKBUF_X1 hold93 (.A(_118_),
    .Z(net93));
 CLKBUF_X1 hold94 (.A(_120_),
    .Z(net94));
 CLKBUF_X1 hold95 (.A(_129_),
    .Z(net95));
 CLKBUF_X1 hold96 (.A(_130_),
    .Z(net96));
 CLKBUF_X1 hold97 (.A(_006_),
    .Z(net97));
 CLKBUF_X1 hold98 (.A(b[1]),
    .Z(net98));
 CLKBUF_X1 hold99 (.A(net33),
    .Z(net99));
 CLKBUF_X1 hold100 (.A(_141_),
    .Z(net100));
 CLKBUF_X1 hold101 (.A(_143_),
    .Z(net101));
 CLKBUF_X1 hold102 (.A(net143),
    .Z(net102));
 CLKBUF_X1 hold103 (.A(_007_),
    .Z(net103));
 CLKBUF_X1 hold104 (.A(b[6]),
    .Z(net104));
 CLKBUF_X1 hold105 (.A(_182_),
    .Z(net105));
 CLKBUF_X1 hold106 (.A(_157_),
    .Z(net106));
 CLKBUF_X1 hold107 (.A(a[3]),
    .Z(net107));
 CLKBUF_X1 hold108 (.A(_189_),
    .Z(net108));
 CLKBUF_X1 hold109 (.A(_190_),
    .Z(net109));
 CLKBUF_X1 hold110 (.A(_097_),
    .Z(net110));
 CLKBUF_X1 hold111 (.A(_098_),
    .Z(net111));
 CLKBUF_X1 hold112 (.A(_099_),
    .Z(net112));
 CLKBUF_X1 hold113 (.A(_004_),
    .Z(net113));
 CLKBUF_X1 hold114 (.A(b[4]),
    .Z(net114));
 CLKBUF_X1 hold115 (.A(_110_),
    .Z(net115));
 CLKBUF_X1 hold116 (.A(_115_),
    .Z(net116));
 CLKBUF_X1 hold117 (.A(net145),
    .Z(net117));
 CLKBUF_X1 hold118 (.A(net118),
    .Z(result[4]));
 CLKBUF_X1 hold119 (.A(net146),
    .Z(net119));
 CLKBUF_X1 hold120 (.A(net120),
    .Z(zero_flag));
 CLKBUF_X1 hold121 (.A(net147),
    .Z(net121));
 CLKBUF_X1 hold122 (.A(net122),
    .Z(result[3]));
 CLKBUF_X1 hold123 (.A(net149),
    .Z(net123));
 CLKBUF_X1 hold124 (.A(net124),
    .Z(result[5]));
 CLKBUF_X1 hold125 (.A(net148),
    .Z(net125));
 CLKBUF_X1 hold126 (.A(net126),
    .Z(result[7]));
 CLKBUF_X1 hold127 (.A(net150),
    .Z(net127));
 CLKBUF_X1 hold128 (.A(net128),
    .Z(result[6]));
 CLKBUF_X1 hold129 (.A(net151),
    .Z(net129));
 CLKBUF_X1 hold130 (.A(net130),
    .Z(result[0]));
 CLKBUF_X1 hold131 (.A(net152),
    .Z(net131));
 CLKBUF_X1 hold132 (.A(net132),
    .Z(result[1]));
 CLKBUF_X1 hold133 (.A(net153),
    .Z(net133));
 CLKBUF_X1 hold134 (.A(net134),
    .Z(result[2]));
 CLKBUF_X1 hold135 (.A(net154),
    .Z(net135));
 CLKBUF_X1 hold136 (.A(net136),
    .Z(overflow_flag));
 CLKBUF_X1 hold137 (.A(opcode[0]),
    .Z(net137));
 CLKBUF_X1 hold138 (.A(a[2]),
    .Z(net138));
 CLKBUF_X1 hold139 (.A(_081_),
    .Z(net139));
 CLKBUF_X1 hold140 (.A(_084_),
    .Z(net140));
 CLKBUF_X1 hold141 (.A(a[5]),
    .Z(net141));
 CLKBUF_X1 hold142 (.A(_214_),
    .Z(net142));
 CLKBUF_X1 hold143 (.A(_144_),
    .Z(net143));
 CLKBUF_X1 hold144 (.A(opcode[3]),
    .Z(net144));
 CLKBUF_X1 hold145 (.A(net55),
    .Z(net145));
 CLKBUF_X1 hold146 (.A(net56),
    .Z(net146));
 CLKBUF_X1 hold147 (.A(net57),
    .Z(net147));
 CLKBUF_X1 hold148 (.A(net59),
    .Z(net148));
 CLKBUF_X1 hold149 (.A(net58),
    .Z(net149));
 CLKBUF_X1 hold150 (.A(net60),
    .Z(net150));
 CLKBUF_X1 hold151 (.A(net61),
    .Z(net151));
 CLKBUF_X1 hold152 (.A(net62),
    .Z(net152));
 CLKBUF_X1 hold153 (.A(net63),
    .Z(net153));
 CLKBUF_X1 hold154 (.A(net64),
    .Z(net154));
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_73 ();
 FILLCELL_X1 FILLER_0_77 ();
 FILLCELL_X32 FILLER_0_79 ();
 FILLCELL_X32 FILLER_0_111 ();
 FILLCELL_X8 FILLER_0_143 ();
 FILLCELL_X4 FILLER_0_151 ();
 FILLCELL_X1 FILLER_0_155 ();
 FILLCELL_X32 FILLER_0_157 ();
 FILLCELL_X32 FILLER_0_189 ();
 FILLCELL_X8 FILLER_0_221 ();
 FILLCELL_X4 FILLER_0_229 ();
 FILLCELL_X1 FILLER_0_233 ();
 FILLCELL_X16 FILLER_0_235 ();
 FILLCELL_X8 FILLER_0_251 ();
 FILLCELL_X2 FILLER_0_259 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X16 FILLER_1_129 ();
 FILLCELL_X8 FILLER_1_145 ();
 FILLCELL_X4 FILLER_1_153 ();
 FILLCELL_X32 FILLER_1_158 ();
 FILLCELL_X32 FILLER_1_190 ();
 FILLCELL_X32 FILLER_1_222 ();
 FILLCELL_X4 FILLER_1_254 ();
 FILLCELL_X2 FILLER_1_258 ();
 FILLCELL_X1 FILLER_1_260 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_73 ();
 FILLCELL_X1 FILLER_2_77 ();
 FILLCELL_X32 FILLER_2_79 ();
 FILLCELL_X32 FILLER_2_111 ();
 FILLCELL_X32 FILLER_2_143 ();
 FILLCELL_X32 FILLER_2_175 ();
 FILLCELL_X16 FILLER_2_207 ();
 FILLCELL_X8 FILLER_2_223 ();
 FILLCELL_X4 FILLER_2_231 ();
 FILLCELL_X16 FILLER_2_236 ();
 FILLCELL_X8 FILLER_2_252 ();
 FILLCELL_X1 FILLER_2_260 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X16 FILLER_3_129 ();
 FILLCELL_X8 FILLER_3_145 ();
 FILLCELL_X4 FILLER_3_153 ();
 FILLCELL_X32 FILLER_3_158 ();
 FILLCELL_X32 FILLER_3_190 ();
 FILLCELL_X32 FILLER_3_222 ();
 FILLCELL_X4 FILLER_3_254 ();
 FILLCELL_X2 FILLER_3_258 ();
 FILLCELL_X1 FILLER_3_260 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X8 FILLER_4_65 ();
 FILLCELL_X4 FILLER_4_73 ();
 FILLCELL_X1 FILLER_4_77 ();
 FILLCELL_X32 FILLER_4_79 ();
 FILLCELL_X32 FILLER_4_111 ();
 FILLCELL_X32 FILLER_4_143 ();
 FILLCELL_X32 FILLER_4_175 ();
 FILLCELL_X16 FILLER_4_207 ();
 FILLCELL_X8 FILLER_4_223 ();
 FILLCELL_X4 FILLER_4_231 ();
 FILLCELL_X16 FILLER_4_236 ();
 FILLCELL_X8 FILLER_4_252 ();
 FILLCELL_X1 FILLER_4_260 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X16 FILLER_5_129 ();
 FILLCELL_X8 FILLER_5_145 ();
 FILLCELL_X4 FILLER_5_153 ();
 FILLCELL_X32 FILLER_5_158 ();
 FILLCELL_X32 FILLER_5_190 ();
 FILLCELL_X32 FILLER_5_222 ();
 FILLCELL_X4 FILLER_5_254 ();
 FILLCELL_X2 FILLER_5_258 ();
 FILLCELL_X1 FILLER_5_260 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X4 FILLER_6_73 ();
 FILLCELL_X1 FILLER_6_77 ();
 FILLCELL_X32 FILLER_6_79 ();
 FILLCELL_X32 FILLER_6_111 ();
 FILLCELL_X32 FILLER_6_143 ();
 FILLCELL_X32 FILLER_6_175 ();
 FILLCELL_X16 FILLER_6_207 ();
 FILLCELL_X8 FILLER_6_223 ();
 FILLCELL_X4 FILLER_6_231 ();
 FILLCELL_X16 FILLER_6_236 ();
 FILLCELL_X8 FILLER_6_252 ();
 FILLCELL_X1 FILLER_6_260 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X16 FILLER_7_129 ();
 FILLCELL_X8 FILLER_7_145 ();
 FILLCELL_X4 FILLER_7_153 ();
 FILLCELL_X32 FILLER_7_158 ();
 FILLCELL_X32 FILLER_7_190 ();
 FILLCELL_X32 FILLER_7_222 ();
 FILLCELL_X4 FILLER_7_254 ();
 FILLCELL_X2 FILLER_7_258 ();
 FILLCELL_X1 FILLER_7_260 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_73 ();
 FILLCELL_X1 FILLER_8_77 ();
 FILLCELL_X32 FILLER_8_79 ();
 FILLCELL_X32 FILLER_8_111 ();
 FILLCELL_X32 FILLER_8_143 ();
 FILLCELL_X32 FILLER_8_175 ();
 FILLCELL_X16 FILLER_8_207 ();
 FILLCELL_X8 FILLER_8_223 ();
 FILLCELL_X4 FILLER_8_231 ();
 FILLCELL_X16 FILLER_8_236 ();
 FILLCELL_X8 FILLER_8_252 ();
 FILLCELL_X1 FILLER_8_260 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X8 FILLER_9_81 ();
 FILLCELL_X4 FILLER_9_89 ();
 FILLCELL_X8 FILLER_9_95 ();
 FILLCELL_X4 FILLER_9_103 ();
 FILLCELL_X1 FILLER_9_107 ();
 FILLCELL_X1 FILLER_9_117 ();
 FILLCELL_X4 FILLER_9_121 ();
 FILLCELL_X16 FILLER_9_127 ();
 FILLCELL_X8 FILLER_9_143 ();
 FILLCELL_X4 FILLER_9_151 ();
 FILLCELL_X2 FILLER_9_155 ();
 FILLCELL_X32 FILLER_9_158 ();
 FILLCELL_X32 FILLER_9_190 ();
 FILLCELL_X32 FILLER_9_222 ();
 FILLCELL_X4 FILLER_9_254 ();
 FILLCELL_X2 FILLER_9_258 ();
 FILLCELL_X1 FILLER_9_260 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_73 ();
 FILLCELL_X1 FILLER_10_77 ();
 FILLCELL_X4 FILLER_10_79 ();
 FILLCELL_X2 FILLER_10_83 ();
 FILLCELL_X4 FILLER_10_104 ();
 FILLCELL_X2 FILLER_10_108 ();
 FILLCELL_X32 FILLER_10_139 ();
 FILLCELL_X32 FILLER_10_171 ();
 FILLCELL_X32 FILLER_10_203 ();
 FILLCELL_X16 FILLER_10_236 ();
 FILLCELL_X8 FILLER_10_252 ();
 FILLCELL_X1 FILLER_10_260 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_33 ();
 FILLCELL_X8 FILLER_11_48 ();
 FILLCELL_X4 FILLER_11_56 ();
 FILLCELL_X4 FILLER_11_62 ();
 FILLCELL_X2 FILLER_11_66 ();
 FILLCELL_X16 FILLER_11_70 ();
 FILLCELL_X8 FILLER_11_86 ();
 FILLCELL_X4 FILLER_11_94 ();
 FILLCELL_X2 FILLER_11_98 ();
 FILLCELL_X1 FILLER_11_100 ();
 FILLCELL_X1 FILLER_11_108 ();
 FILLCELL_X16 FILLER_11_139 ();
 FILLCELL_X2 FILLER_11_155 ();
 FILLCELL_X32 FILLER_11_158 ();
 FILLCELL_X32 FILLER_11_190 ();
 FILLCELL_X32 FILLER_11_222 ();
 FILLCELL_X4 FILLER_11_254 ();
 FILLCELL_X2 FILLER_11_258 ();
 FILLCELL_X1 FILLER_11_260 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_17 ();
 FILLCELL_X4 FILLER_12_25 ();
 FILLCELL_X2 FILLER_12_29 ();
 FILLCELL_X1 FILLER_12_31 ();
 FILLCELL_X2 FILLER_12_59 ();
 FILLCELL_X4 FILLER_12_64 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X2 FILLER_12_113 ();
 FILLCELL_X1 FILLER_12_115 ();
 FILLCELL_X1 FILLER_12_124 ();
 FILLCELL_X8 FILLER_12_128 ();
 FILLCELL_X2 FILLER_12_136 ();
 FILLCELL_X1 FILLER_12_138 ();
 FILLCELL_X32 FILLER_12_153 ();
 FILLCELL_X32 FILLER_12_185 ();
 FILLCELL_X16 FILLER_12_217 ();
 FILLCELL_X2 FILLER_12_233 ();
 FILLCELL_X16 FILLER_12_236 ();
 FILLCELL_X8 FILLER_12_252 ();
 FILLCELL_X1 FILLER_12_260 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_9 ();
 FILLCELL_X4 FILLER_13_16 ();
 FILLCELL_X2 FILLER_13_20 ();
 FILLCELL_X1 FILLER_13_22 ();
 FILLCELL_X1 FILLER_13_33 ();
 FILLCELL_X1 FILLER_13_44 ();
 FILLCELL_X16 FILLER_13_50 ();
 FILLCELL_X2 FILLER_13_66 ();
 FILLCELL_X1 FILLER_13_68 ();
 FILLCELL_X8 FILLER_13_72 ();
 FILLCELL_X2 FILLER_13_93 ();
 FILLCELL_X1 FILLER_13_95 ();
 FILLCELL_X8 FILLER_13_100 ();
 FILLCELL_X4 FILLER_13_108 ();
 FILLCELL_X1 FILLER_13_116 ();
 FILLCELL_X1 FILLER_13_126 ();
 FILLCELL_X1 FILLER_13_134 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X4 FILLER_13_257 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_9 ();
 FILLCELL_X2 FILLER_14_13 ();
 FILLCELL_X1 FILLER_14_15 ();
 FILLCELL_X8 FILLER_14_27 ();
 FILLCELL_X2 FILLER_14_35 ();
 FILLCELL_X1 FILLER_14_45 ();
 FILLCELL_X2 FILLER_14_57 ();
 FILLCELL_X8 FILLER_14_66 ();
 FILLCELL_X4 FILLER_14_74 ();
 FILLCELL_X2 FILLER_14_105 ();
 FILLCELL_X1 FILLER_14_112 ();
 FILLCELL_X2 FILLER_14_121 ();
 FILLCELL_X1 FILLER_14_123 ();
 FILLCELL_X16 FILLER_14_130 ();
 FILLCELL_X32 FILLER_14_155 ();
 FILLCELL_X32 FILLER_14_187 ();
 FILLCELL_X16 FILLER_14_219 ();
 FILLCELL_X16 FILLER_14_236 ();
 FILLCELL_X8 FILLER_14_252 ();
 FILLCELL_X1 FILLER_14_260 ();
 FILLCELL_X1 FILLER_15_4 ();
 FILLCELL_X8 FILLER_15_49 ();
 FILLCELL_X2 FILLER_15_57 ();
 FILLCELL_X8 FILLER_15_75 ();
 FILLCELL_X2 FILLER_15_83 ();
 FILLCELL_X1 FILLER_15_85 ();
 FILLCELL_X2 FILLER_15_93 ();
 FILLCELL_X4 FILLER_15_100 ();
 FILLCELL_X2 FILLER_15_104 ();
 FILLCELL_X1 FILLER_15_106 ();
 FILLCELL_X4 FILLER_15_125 ();
 FILLCELL_X2 FILLER_15_129 ();
 FILLCELL_X4 FILLER_15_136 ();
 FILLCELL_X2 FILLER_15_140 ();
 FILLCELL_X1 FILLER_15_142 ();
 FILLCELL_X4 FILLER_15_153 ();
 FILLCELL_X8 FILLER_15_165 ();
 FILLCELL_X2 FILLER_15_173 ();
 FILLCELL_X1 FILLER_15_175 ();
 FILLCELL_X32 FILLER_15_195 ();
 FILLCELL_X32 FILLER_15_227 ();
 FILLCELL_X2 FILLER_15_259 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_17 ();
 FILLCELL_X2 FILLER_16_22 ();
 FILLCELL_X4 FILLER_16_49 ();
 FILLCELL_X2 FILLER_16_53 ();
 FILLCELL_X4 FILLER_16_58 ();
 FILLCELL_X1 FILLER_16_62 ();
 FILLCELL_X8 FILLER_16_68 ();
 FILLCELL_X2 FILLER_16_76 ();
 FILLCELL_X2 FILLER_16_79 ();
 FILLCELL_X1 FILLER_16_86 ();
 FILLCELL_X2 FILLER_16_91 ();
 FILLCELL_X16 FILLER_16_110 ();
 FILLCELL_X2 FILLER_16_126 ();
 FILLCELL_X1 FILLER_16_128 ();
 FILLCELL_X8 FILLER_16_134 ();
 FILLCELL_X2 FILLER_16_142 ();
 FILLCELL_X4 FILLER_16_153 ();
 FILLCELL_X4 FILLER_16_163 ();
 FILLCELL_X2 FILLER_16_167 ();
 FILLCELL_X1 FILLER_16_169 ();
 FILLCELL_X2 FILLER_16_177 ();
 FILLCELL_X8 FILLER_16_198 ();
 FILLCELL_X2 FILLER_16_206 ();
 FILLCELL_X1 FILLER_16_208 ();
 FILLCELL_X8 FILLER_16_212 ();
 FILLCELL_X4 FILLER_16_220 ();
 FILLCELL_X8 FILLER_16_227 ();
 FILLCELL_X16 FILLER_16_236 ();
 FILLCELL_X4 FILLER_16_252 ();
 FILLCELL_X2 FILLER_16_259 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_9 ();
 FILLCELL_X2 FILLER_17_17 ();
 FILLCELL_X8 FILLER_17_25 ();
 FILLCELL_X2 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_38 ();
 FILLCELL_X1 FILLER_17_48 ();
 FILLCELL_X2 FILLER_17_55 ();
 FILLCELL_X1 FILLER_17_57 ();
 FILLCELL_X2 FILLER_17_63 ();
 FILLCELL_X1 FILLER_17_65 ();
 FILLCELL_X4 FILLER_17_74 ();
 FILLCELL_X2 FILLER_17_78 ();
 FILLCELL_X1 FILLER_17_80 ();
 FILLCELL_X1 FILLER_17_87 ();
 FILLCELL_X4 FILLER_17_114 ();
 FILLCELL_X1 FILLER_17_118 ();
 FILLCELL_X2 FILLER_17_126 ();
 FILLCELL_X2 FILLER_17_138 ();
 FILLCELL_X1 FILLER_17_153 ();
 FILLCELL_X1 FILLER_17_158 ();
 FILLCELL_X16 FILLER_17_193 ();
 FILLCELL_X2 FILLER_17_209 ();
 FILLCELL_X1 FILLER_17_211 ();
 FILLCELL_X8 FILLER_17_215 ();
 FILLCELL_X4 FILLER_17_223 ();
 FILLCELL_X16 FILLER_17_230 ();
 FILLCELL_X1 FILLER_17_246 ();
 FILLCELL_X2 FILLER_17_256 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_27 ();
 FILLCELL_X2 FILLER_18_36 ();
 FILLCELL_X32 FILLER_18_42 ();
 FILLCELL_X4 FILLER_18_74 ();
 FILLCELL_X16 FILLER_18_79 ();
 FILLCELL_X1 FILLER_18_109 ();
 FILLCELL_X8 FILLER_18_113 ();
 FILLCELL_X4 FILLER_18_121 ();
 FILLCELL_X2 FILLER_18_125 ();
 FILLCELL_X1 FILLER_18_129 ();
 FILLCELL_X1 FILLER_18_139 ();
 FILLCELL_X2 FILLER_18_142 ();
 FILLCELL_X8 FILLER_18_147 ();
 FILLCELL_X4 FILLER_18_155 ();
 FILLCELL_X2 FILLER_18_159 ();
 FILLCELL_X1 FILLER_18_161 ();
 FILLCELL_X4 FILLER_18_165 ();
 FILLCELL_X2 FILLER_18_169 ();
 FILLCELL_X1 FILLER_18_171 ();
 FILLCELL_X8 FILLER_18_177 ();
 FILLCELL_X4 FILLER_18_185 ();
 FILLCELL_X2 FILLER_18_189 ();
 FILLCELL_X1 FILLER_18_191 ();
 FILLCELL_X8 FILLER_18_197 ();
 FILLCELL_X2 FILLER_18_205 ();
 FILLCELL_X1 FILLER_18_207 ();
 FILLCELL_X8 FILLER_18_211 ();
 FILLCELL_X4 FILLER_18_219 ();
 FILLCELL_X8 FILLER_18_226 ();
 FILLCELL_X1 FILLER_18_234 ();
 FILLCELL_X8 FILLER_18_236 ();
 FILLCELL_X2 FILLER_18_244 ();
 FILLCELL_X16 FILLER_19_4 ();
 FILLCELL_X8 FILLER_19_20 ();
 FILLCELL_X4 FILLER_19_28 ();
 FILLCELL_X2 FILLER_19_32 ();
 FILLCELL_X1 FILLER_19_37 ();
 FILLCELL_X4 FILLER_19_41 ();
 FILLCELL_X2 FILLER_19_45 ();
 FILLCELL_X4 FILLER_19_50 ();
 FILLCELL_X1 FILLER_19_54 ();
 FILLCELL_X16 FILLER_19_74 ();
 FILLCELL_X8 FILLER_19_90 ();
 FILLCELL_X4 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_102 ();
 FILLCELL_X2 FILLER_19_107 ();
 FILLCELL_X1 FILLER_19_109 ();
 FILLCELL_X2 FILLER_19_116 ();
 FILLCELL_X8 FILLER_19_130 ();
 FILLCELL_X2 FILLER_19_138 ();
 FILLCELL_X4 FILLER_19_143 ();
 FILLCELL_X2 FILLER_19_147 ();
 FILLCELL_X1 FILLER_19_156 ();
 FILLCELL_X4 FILLER_19_158 ();
 FILLCELL_X2 FILLER_19_162 ();
 FILLCELL_X1 FILLER_19_169 ();
 FILLCELL_X2 FILLER_19_177 ();
 FILLCELL_X1 FILLER_19_179 ();
 FILLCELL_X16 FILLER_19_199 ();
 FILLCELL_X8 FILLER_19_215 ();
 FILLCELL_X4 FILLER_19_223 ();
 FILLCELL_X16 FILLER_19_230 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_24 ();
 FILLCELL_X1 FILLER_20_26 ();
 FILLCELL_X2 FILLER_20_44 ();
 FILLCELL_X8 FILLER_20_59 ();
 FILLCELL_X2 FILLER_20_67 ();
 FILLCELL_X1 FILLER_20_74 ();
 FILLCELL_X2 FILLER_20_79 ();
 FILLCELL_X2 FILLER_20_104 ();
 FILLCELL_X1 FILLER_20_106 ();
 FILLCELL_X4 FILLER_20_125 ();
 FILLCELL_X1 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_132 ();
 FILLCELL_X2 FILLER_20_140 ();
 FILLCELL_X1 FILLER_20_142 ();
 FILLCELL_X1 FILLER_20_152 ();
 FILLCELL_X2 FILLER_20_175 ();
 FILLCELL_X8 FILLER_20_202 ();
 FILLCELL_X4 FILLER_20_210 ();
 FILLCELL_X1 FILLER_20_214 ();
 FILLCELL_X8 FILLER_20_221 ();
 FILLCELL_X1 FILLER_20_229 ();
 FILLCELL_X2 FILLER_20_233 ();
 FILLCELL_X8 FILLER_20_236 ();
 FILLCELL_X4 FILLER_20_244 ();
 FILLCELL_X1 FILLER_20_251 ();
 FILLCELL_X1 FILLER_20_255 ();
 FILLCELL_X2 FILLER_20_259 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_9 ();
 FILLCELL_X4 FILLER_21_21 ();
 FILLCELL_X1 FILLER_21_25 ();
 FILLCELL_X4 FILLER_21_29 ();
 FILLCELL_X2 FILLER_21_33 ();
 FILLCELL_X1 FILLER_21_35 ();
 FILLCELL_X8 FILLER_21_40 ();
 FILLCELL_X4 FILLER_21_48 ();
 FILLCELL_X2 FILLER_21_52 ();
 FILLCELL_X4 FILLER_21_58 ();
 FILLCELL_X1 FILLER_21_87 ();
 FILLCELL_X4 FILLER_21_94 ();
 FILLCELL_X1 FILLER_21_98 ();
 FILLCELL_X16 FILLER_21_111 ();
 FILLCELL_X8 FILLER_21_129 ();
 FILLCELL_X1 FILLER_21_137 ();
 FILLCELL_X2 FILLER_21_155 ();
 FILLCELL_X4 FILLER_21_158 ();
 FILLCELL_X2 FILLER_21_162 ();
 FILLCELL_X1 FILLER_21_164 ();
 FILLCELL_X2 FILLER_21_169 ();
 FILLCELL_X8 FILLER_21_198 ();
 FILLCELL_X4 FILLER_21_206 ();
 FILLCELL_X2 FILLER_21_210 ();
 FILLCELL_X4 FILLER_21_215 ();
 FILLCELL_X2 FILLER_21_219 ();
 FILLCELL_X2 FILLER_21_224 ();
 FILLCELL_X1 FILLER_21_226 ();
 FILLCELL_X8 FILLER_21_230 ();
 FILLCELL_X4 FILLER_21_238 ();
 FILLCELL_X1 FILLER_21_242 ();
 FILLCELL_X8 FILLER_21_249 ();
 FILLCELL_X4 FILLER_21_257 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_23 ();
 FILLCELL_X2 FILLER_22_27 ();
 FILLCELL_X8 FILLER_22_32 ();
 FILLCELL_X4 FILLER_22_40 ();
 FILLCELL_X1 FILLER_22_44 ();
 FILLCELL_X16 FILLER_22_48 ();
 FILLCELL_X4 FILLER_22_68 ();
 FILLCELL_X2 FILLER_22_75 ();
 FILLCELL_X1 FILLER_22_77 ();
 FILLCELL_X2 FILLER_22_79 ();
 FILLCELL_X1 FILLER_22_81 ();
 FILLCELL_X8 FILLER_22_86 ();
 FILLCELL_X4 FILLER_22_94 ();
 FILLCELL_X4 FILLER_22_105 ();
 FILLCELL_X4 FILLER_22_113 ();
 FILLCELL_X2 FILLER_22_117 ();
 FILLCELL_X1 FILLER_22_119 ();
 FILLCELL_X8 FILLER_22_143 ();
 FILLCELL_X1 FILLER_22_166 ();
 FILLCELL_X1 FILLER_22_170 ();
 FILLCELL_X8 FILLER_22_193 ();
 FILLCELL_X4 FILLER_22_201 ();
 FILLCELL_X4 FILLER_22_208 ();
 FILLCELL_X2 FILLER_22_212 ();
 FILLCELL_X1 FILLER_22_214 ();
 FILLCELL_X16 FILLER_22_218 ();
 FILLCELL_X1 FILLER_22_234 ();
 FILLCELL_X16 FILLER_22_236 ();
 FILLCELL_X8 FILLER_22_252 ();
 FILLCELL_X1 FILLER_22_260 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_17 ();
 FILLCELL_X4 FILLER_23_25 ();
 FILLCELL_X2 FILLER_23_29 ();
 FILLCELL_X1 FILLER_23_31 ();
 FILLCELL_X2 FILLER_23_36 ();
 FILLCELL_X1 FILLER_23_38 ();
 FILLCELL_X8 FILLER_23_58 ();
 FILLCELL_X4 FILLER_23_66 ();
 FILLCELL_X4 FILLER_23_76 ();
 FILLCELL_X2 FILLER_23_90 ();
 FILLCELL_X4 FILLER_23_96 ();
 FILLCELL_X1 FILLER_23_100 ();
 FILLCELL_X2 FILLER_23_111 ();
 FILLCELL_X1 FILLER_23_113 ();
 FILLCELL_X2 FILLER_23_117 ();
 FILLCELL_X16 FILLER_23_130 ();
 FILLCELL_X4 FILLER_23_146 ();
 FILLCELL_X1 FILLER_23_150 ();
 FILLCELL_X2 FILLER_23_155 ();
 FILLCELL_X2 FILLER_23_162 ();
 FILLCELL_X16 FILLER_23_183 ();
 FILLCELL_X4 FILLER_23_202 ();
 FILLCELL_X2 FILLER_23_206 ();
 FILLCELL_X32 FILLER_23_214 ();
 FILLCELL_X8 FILLER_23_246 ();
 FILLCELL_X4 FILLER_23_254 ();
 FILLCELL_X2 FILLER_23_258 ();
 FILLCELL_X1 FILLER_23_260 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X4 FILLER_24_17 ();
 FILLCELL_X2 FILLER_24_21 ();
 FILLCELL_X1 FILLER_24_28 ();
 FILLCELL_X1 FILLER_24_38 ();
 FILLCELL_X4 FILLER_24_52 ();
 FILLCELL_X1 FILLER_24_56 ();
 FILLCELL_X2 FILLER_24_63 ();
 FILLCELL_X16 FILLER_24_125 ();
 FILLCELL_X8 FILLER_24_141 ();
 FILLCELL_X2 FILLER_24_149 ();
 FILLCELL_X16 FILLER_24_173 ();
 FILLCELL_X1 FILLER_24_189 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X8 FILLER_24_225 ();
 FILLCELL_X2 FILLER_24_233 ();
 FILLCELL_X16 FILLER_24_236 ();
 FILLCELL_X8 FILLER_24_252 ();
 FILLCELL_X1 FILLER_24_260 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_33 ();
 FILLCELL_X2 FILLER_25_37 ();
 FILLCELL_X1 FILLER_25_39 ();
 FILLCELL_X8 FILLER_25_50 ();
 FILLCELL_X4 FILLER_25_58 ();
 FILLCELL_X2 FILLER_25_62 ();
 FILLCELL_X1 FILLER_25_64 ();
 FILLCELL_X2 FILLER_25_74 ();
 FILLCELL_X8 FILLER_25_95 ();
 FILLCELL_X32 FILLER_25_105 ();
 FILLCELL_X16 FILLER_25_137 ();
 FILLCELL_X4 FILLER_25_153 ();
 FILLCELL_X8 FILLER_25_182 ();
 FILLCELL_X4 FILLER_25_190 ();
 FILLCELL_X32 FILLER_25_197 ();
 FILLCELL_X32 FILLER_25_229 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X16 FILLER_26_33 ();
 FILLCELL_X8 FILLER_26_49 ();
 FILLCELL_X4 FILLER_26_57 ();
 FILLCELL_X1 FILLER_26_61 ();
 FILLCELL_X4 FILLER_26_71 ();
 FILLCELL_X2 FILLER_26_75 ();
 FILLCELL_X1 FILLER_26_77 ();
 FILLCELL_X32 FILLER_26_82 ();
 FILLCELL_X32 FILLER_26_114 ();
 FILLCELL_X16 FILLER_26_146 ();
 FILLCELL_X4 FILLER_26_165 ();
 FILLCELL_X32 FILLER_26_173 ();
 FILLCELL_X16 FILLER_26_205 ();
 FILLCELL_X8 FILLER_26_221 ();
 FILLCELL_X4 FILLER_26_229 ();
 FILLCELL_X2 FILLER_26_233 ();
 FILLCELL_X16 FILLER_26_236 ();
 FILLCELL_X8 FILLER_26_252 ();
 FILLCELL_X1 FILLER_26_260 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X16 FILLER_27_33 ();
 FILLCELL_X8 FILLER_27_49 ();
 FILLCELL_X4 FILLER_27_57 ();
 FILLCELL_X2 FILLER_27_61 ();
 FILLCELL_X32 FILLER_27_74 ();
 FILLCELL_X32 FILLER_27_106 ();
 FILLCELL_X16 FILLER_27_138 ();
 FILLCELL_X2 FILLER_27_154 ();
 FILLCELL_X1 FILLER_27_156 ();
 FILLCELL_X32 FILLER_27_158 ();
 FILLCELL_X32 FILLER_27_190 ();
 FILLCELL_X32 FILLER_27_222 ();
 FILLCELL_X4 FILLER_27_254 ();
 FILLCELL_X2 FILLER_27_258 ();
 FILLCELL_X1 FILLER_27_260 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X8 FILLER_28_65 ();
 FILLCELL_X4 FILLER_28_73 ();
 FILLCELL_X1 FILLER_28_77 ();
 FILLCELL_X32 FILLER_28_79 ();
 FILLCELL_X32 FILLER_28_111 ();
 FILLCELL_X32 FILLER_28_143 ();
 FILLCELL_X32 FILLER_28_175 ();
 FILLCELL_X16 FILLER_28_207 ();
 FILLCELL_X8 FILLER_28_223 ();
 FILLCELL_X4 FILLER_28_231 ();
 FILLCELL_X16 FILLER_28_236 ();
 FILLCELL_X8 FILLER_28_252 ();
 FILLCELL_X1 FILLER_28_260 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X16 FILLER_29_129 ();
 FILLCELL_X8 FILLER_29_145 ();
 FILLCELL_X4 FILLER_29_153 ();
 FILLCELL_X32 FILLER_29_158 ();
 FILLCELL_X32 FILLER_29_190 ();
 FILLCELL_X32 FILLER_29_222 ();
 FILLCELL_X4 FILLER_29_254 ();
 FILLCELL_X2 FILLER_29_258 ();
 FILLCELL_X1 FILLER_29_260 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X8 FILLER_30_65 ();
 FILLCELL_X4 FILLER_30_73 ();
 FILLCELL_X1 FILLER_30_77 ();
 FILLCELL_X32 FILLER_30_79 ();
 FILLCELL_X32 FILLER_30_111 ();
 FILLCELL_X32 FILLER_30_143 ();
 FILLCELL_X32 FILLER_30_175 ();
 FILLCELL_X16 FILLER_30_207 ();
 FILLCELL_X8 FILLER_30_223 ();
 FILLCELL_X4 FILLER_30_231 ();
 FILLCELL_X16 FILLER_30_236 ();
 FILLCELL_X8 FILLER_30_252 ();
 FILLCELL_X1 FILLER_30_260 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X16 FILLER_31_129 ();
 FILLCELL_X8 FILLER_31_145 ();
 FILLCELL_X4 FILLER_31_153 ();
 FILLCELL_X32 FILLER_31_158 ();
 FILLCELL_X32 FILLER_31_190 ();
 FILLCELL_X32 FILLER_31_222 ();
 FILLCELL_X4 FILLER_31_254 ();
 FILLCELL_X2 FILLER_31_258 ();
 FILLCELL_X1 FILLER_31_260 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X8 FILLER_32_65 ();
 FILLCELL_X4 FILLER_32_73 ();
 FILLCELL_X1 FILLER_32_77 ();
 FILLCELL_X32 FILLER_32_79 ();
 FILLCELL_X32 FILLER_32_111 ();
 FILLCELL_X32 FILLER_32_143 ();
 FILLCELL_X32 FILLER_32_175 ();
 FILLCELL_X16 FILLER_32_207 ();
 FILLCELL_X8 FILLER_32_223 ();
 FILLCELL_X4 FILLER_32_231 ();
 FILLCELL_X16 FILLER_32_236 ();
 FILLCELL_X8 FILLER_32_252 ();
 FILLCELL_X1 FILLER_32_260 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X8 FILLER_33_65 ();
 FILLCELL_X4 FILLER_33_73 ();
 FILLCELL_X1 FILLER_33_77 ();
 FILLCELL_X8 FILLER_33_79 ();
 FILLCELL_X4 FILLER_33_87 ();
 FILLCELL_X2 FILLER_33_91 ();
 FILLCELL_X1 FILLER_33_93 ();
 FILLCELL_X8 FILLER_33_103 ();
 FILLCELL_X1 FILLER_33_111 ();
 FILLCELL_X32 FILLER_33_115 ();
 FILLCELL_X8 FILLER_33_147 ();
 FILLCELL_X1 FILLER_33_155 ();
 FILLCELL_X32 FILLER_33_157 ();
 FILLCELL_X32 FILLER_33_189 ();
 FILLCELL_X8 FILLER_33_221 ();
 FILLCELL_X4 FILLER_33_229 ();
 FILLCELL_X1 FILLER_33_233 ();
 FILLCELL_X16 FILLER_33_235 ();
 FILLCELL_X8 FILLER_33_251 ();
 FILLCELL_X2 FILLER_33_259 ();
endmodule
